<?xml version="1.0" encoding="UTF-8"?>
<svg version="1.1" xmlns="http://www.w3.org/2000/svg" width="1024" height="1024">
<path d="M0 0 C337.92 0 675.84 0 1024 0 C1024 337.92 1024 675.84 1024 1024 C686.08 1024 348.16 1024 0 1024 C0 686.08 0 348.16 0 0 Z " fill="#F9F9F9" transform="translate(0,0)"/>
<path d="M0 0 C266.31 0 532.62 0 807 0 C807 232.65 807 465.3 807 705 C789.18 705 771.36 705 753 705 C753 722.49 753 739.98 753 758 C735.18 758 717.36 758 699 758 C699 775.49 699 792.98 699 811 C681.51 811 664.02 811 646 811 C646 828.49 646 845.98 646 864 C632.9134375 864.0309375 632.9134375 864.0309375 619.5625 864.0625 C616.80463135 864.071604 614.0467627 864.08070801 611.20532227 864.09008789 C609.03401742 864.09300684 606.86271204 864.09555545 604.69140625 864.09765625 C603.55215698 864.10277222 602.41290771 864.10788818 601.23913574 864.11315918 C600.16321167 864.11328003 599.0872876 864.11340088 597.97875977 864.11352539 C596.56978172 864.11685631 596.56978172 864.11685631 595.13233948 864.12025452 C593 864 593 864 592 863 C591.90659566 861.37325222 591.88254829 859.74245949 591.88647461 858.11303711 C591.88665588 856.5296051 591.88665588 856.5296051 591.88684082 854.91418457 C591.89451477 853.23769836 591.89451477 853.23769836 591.90234375 851.52734375 C591.90335083 850.50612427 591.90435791 849.48490479 591.90539551 848.43273926 C591.91064585 844.60098149 591.92460697 840.76923967 591.9375 836.9375 C591.958125 828.378125 591.97875 819.81875 592 811 C574.18 811 556.36 811 538 811 C537.67 793.51 537.34 776.02 537 758 C564.225 757.505 564.225 757.505 592 757 C591.96040949 740.96409456 591.96040949 740.96409456 591.90991211 724.92822266 C591.90699254 722.92350314 591.90444408 720.91878304 591.90234375 718.9140625 C591.89722778 717.86629639 591.89211182 716.81853027 591.88684082 715.73901367 C591.88671997 714.74442139 591.88659912 713.7498291 591.88647461 712.72509766 C591.884254 711.85905914 591.88203339 710.99302063 591.87974548 710.10073853 C592 708 592 708 593 706 C610.68978255 704.88442813 628.27711691 704.92458348 646 705 C646 687.84 646 670.68 646 653 C663.49 653 680.98 653 699 653 C699 635.51 699 618.02 699 600 C681.51 600 664.02 600 646 600 C645.9690625 587.1609375 645.9690625 587.1609375 645.9375 574.0625 C645.928396 571.35683838 645.91929199 568.65117676 645.90991211 565.86352539 C645.90699315 563.73323618 645.90444455 561.60294642 645.90234375 559.47265625 C645.89722778 558.35499878 645.89211182 557.23734131 645.88684082 556.08581543 C645.88671997 555.03019409 645.88659912 553.97457275 645.88647461 552.88696289 C645.884254 551.96540909 645.88203339 551.04385529 645.87974548 550.09437561 C646 548 646 548 647 547 C648.62674778 546.90659566 650.25754051 546.88254829 651.88696289 546.88647461 C653.4703949 546.88665588 653.4703949 546.88665588 655.08581543 546.88684082 C656.76230164 546.89451477 656.76230164 546.89451477 658.47265625 546.90234375 C660.00448547 546.90385437 660.00448547 546.90385437 661.56726074 546.90539551 C665.39901851 546.91064585 669.23076033 546.92460697 673.0625 546.9375 C681.621875 546.958125 690.18125 546.97875 699 547 C699 529.84 699 512.68 699 495 C681.51 495 664.02 495 646 495 C646 512.16 646 529.32 646 547 C643.51644959 548.24177521 641.86892378 548.12036681 639.09130859 548.11352539 C638.07040131 548.11344986 637.04949402 548.11337433 635.99765015 548.11329651 C634.33978989 548.10555458 634.33978989 548.10555458 632.6484375 548.09765625 C631.5192691 548.0962413 630.39010071 548.09482635 629.22671509 548.09336853 C625.60945012 548.08775744 621.99224636 548.07520303 618.375 548.0625 C615.92708423 548.05748643 613.47916748 548.05292328 611.03125 548.04882812 C605.02081234 548.0377844 599.01041054 548.02103544 593 548 C593.00333092 548.82232872 593.00333092 548.82232872 593.00672913 549.66127014 C593.02892226 555.38802435 593.04396499 561.11476626 593.05493164 566.84155273 C593.05994778 568.97632341 593.06676224 571.11109067 593.07543945 573.24584961 C593.08762435 576.32146042 593.09325562 579.39702563 593.09765625 582.47265625 C593.10281754 583.42084732 593.10797882 584.36903839 593.11329651 585.34596252 C593.11337204 586.24636765 593.11344757 587.14677277 593.11352539 588.07446289 C593.115746 588.85833878 593.11796661 589.64221466 593.12025452 590.44984436 C592.9692781 593.65149841 592.4532854 596.82700222 592 600 C574.51 600 557.02 600 539 600 C538.13520548 544.9414158 538.13520548 544.9414158 544.27685547 525.48266602 C560.28209595 470.53422225 544.5806975 405.37352229 518.109375 356.48828125 C508.78421483 339.7480392 497.28336475 324.44713465 484.24609375 310.43359375 C482.36544087 308.39594724 480.58355404 306.31907394 478.8125 304.1875 C452.66592445 274.13752573 412.41509735 248.53865503 374 238 C374.66 237.67 375.32 237.34 376 237 C377.190189 232.93924972 377.12079049 228.93769286 377.11352539 224.73120117 C377.11374443 223.66209 377.11374443 223.66209 377.1139679 222.57138062 C377.11327432 220.2285451 377.105508 217.88579028 377.09765625 215.54296875 C377.0957901 213.91343733 377.09436713 212.28390535 377.09336853 210.65437317 C377.08955888 206.37511636 377.07974188 202.09589374 377.06866455 197.81665039 C377.05661384 192.67708289 377.0520408 187.53750393 377.04621124 182.39792633 C377.03652927 174.59859381 377.01736187 166.79933624 377 159 C359.18 159 341.36 159 323 159 C323 176.16 323 193.32 323 211 C305.18 211 287.36 211 269 211 C269 193.84 269 176.68 269 159 C251.51 159.33 234.02 159.66 216 160 C215.67 176.83 215.34 193.66 215 211 C197.51 211 180.02 211 162 211 C162 193.84 162 176.68 162 159 C179.49 159 196.98 159 215 159 C214.9603903 141.93174701 214.9603903 141.93174701 214.90991211 124.86352539 C214.90699315 122.73323618 214.90444455 120.60294642 214.90234375 118.47265625 C214.89722778 117.35499878 214.89211182 116.23734131 214.88684082 115.08581543 C214.88665955 113.50238342 214.88665955 113.50238342 214.88647461 111.88696289 C214.884254 110.96540909 214.88203339 110.04385529 214.87974548 109.09437561 C215 107 215 107 216 106 C217.65738443 105.90653085 219.31874644 105.88255023 220.97875977 105.88647461 C222.05468384 105.88659546 223.13060791 105.88671631 224.23913574 105.88684082 C225.37838501 105.89195679 226.51763428 105.89707275 227.69140625 105.90234375 C229.25272278 105.90385437 229.25272278 105.90385437 230.84558105 105.90539551 C234.75123184 105.91064599 238.65686697 105.92460711 242.5625 105.9375 C251.286875 105.958125 260.01125 105.97875 269 106 C269 88.51 269 71.02 269 53 C251.18 53 233.36 53 215 53 C215 70.49 215 87.98 215 106 C197.51 106 180.02 106 162 106 C162 88.51 162 71.02 162 53 C143.85 53 125.7 53 107 53 C107 70.49 107 87.98 107 106 C89.51 106 72.02 106 54 106 C54 88.51 54 71.02 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FBFBFB" transform="translate(217,0)"/>
<path d="M0 0 C0.92141785 -0.00701431 1.84283569 -0.01402863 2.79217529 -0.02125549 C5.75603156 -0.03869159 8.71968804 -0.04510954 11.68359375 -0.046875 C13.20199356 -0.04788712 13.20199356 -0.04788712 14.75106812 -0.04891968 C29.7752844 -0.03298984 44.31596387 0.44362914 59.12109375 3.203125 C60.08063965 3.36941406 61.04018555 3.53570312 62.02880859 3.70703125 C84.02343127 7.56010384 105.06616841 14.38909993 125.12109375 24.203125 C126.01151367 24.63608887 126.90193359 25.06905273 127.81933594 25.51513672 C186.52710837 54.34717607 235.36620413 106.64948816 257.05859375 168.765625 C258.11740692 171.90010402 259.13367147 175.04548209 260.12109375 178.203125 C260.32814941 178.86135254 260.53520508 179.51958008 260.74853516 180.19775391 C264.32069212 191.714725 266.70564405 203.45778078 268.74609375 215.328125 C268.86927979 216.03163086 268.99246582 216.73513672 269.11938477 217.45996094 C275.30584129 254.68985964 271.29642037 296.86104155 258.12109375 332.203125 C257.79157715 333.09854004 257.46206055 333.99395508 257.12255859 334.91650391 C248.96730591 356.8174475 239.02469021 377.37167156 225.12109375 396.203125 C224.33001305 397.30026525 223.53962365 398.39790438 222.75 399.49609375 C217.91405607 406.10884897 212.67752814 412.19172125 207.12109375 418.203125 C205.66179636 419.8481036 204.20347065 421.49394469 202.74609375 423.140625 C194.49206878 432.28310405 185.85157861 440.64607322 176.12109375 448.203125 C175.5585791 448.64736816 174.99606445 449.09161133 174.41650391 449.54931641 C145.97735913 471.94869685 113.26113681 488.11313987 78.18676758 497.17700195 C75.58718686 497.85019672 75.58718686 497.85019672 72.12109375 499.203125 C70.97422075 501.2000588 70.97422075 501.2000588 70.12109375 503.203125 C65.92963909 505.13300341 60.59575896 504.24734434 56.05273438 504.1640625 C52.16043789 504.12028784 48.98676122 504.42999151 45.12109375 505.203125 C44.79109375 514.443125 44.46109375 523.683125 44.12109375 533.203125 C45.11109375 533.533125 46.10109375 533.863125 47.12109375 534.203125 C46.46109375 534.533125 45.80109375 534.863125 45.12109375 535.203125 C44.79109375 552.033125 44.46109375 568.863125 44.12109375 586.203125 C26.63109375 586.533125 9.14109375 586.863125 -8.87890625 587.203125 C-9.20890625 604.363125 -9.53890625 621.523125 -9.87890625 639.203125 C-45.18890625 639.203125 -80.49890625 639.203125 -116.87890625 639.203125 C-116.87890625 622.043125 -116.87890625 604.883125 -116.87890625 587.203125 C-134.69890625 586.873125 -152.51890625 586.543125 -170.87890625 586.203125 C-170.89953125 577.64375 -170.92015625 569.084375 -170.94140625 560.265625 C-170.95051025 557.55996338 -170.95961426 554.85430176 -170.96899414 552.06665039 C-170.9719131 549.93636118 -170.9744617 547.80607142 -170.9765625 545.67578125 C-170.98167847 544.55812378 -170.98679443 543.44046631 -170.99206543 542.28894043 C-170.9922467 540.70550842 -170.9922467 540.70550842 -170.99243164 539.09008789 C-170.99465225 538.16853409 -170.99687286 537.24698029 -170.99916077 536.29750061 C-170.87890625 534.203125 -170.87890625 534.203125 -169.87890625 533.203125 C-168.22152182 533.10965585 -166.56015981 533.08567523 -164.90014648 533.08959961 C-163.83912216 533.08967514 -162.77809784 533.08975067 -161.68492126 533.08982849 C-160.53077225 533.09498978 -159.37662323 533.10015106 -158.1875 533.10546875 C-157.01252457 533.1068837 -155.83754913 533.10829865 -154.62696838 533.10975647 C-150.85675561 533.11537508 -147.08660121 533.12793074 -143.31640625 533.140625 C-140.76757898 533.1456376 -138.21875078 533.15020092 -135.66992188 533.15429688 C-129.40620916 533.16450169 -123.14262341 533.18407348 -116.87890625 533.203125 C-116.87890625 516.043125 -116.87890625 498.883125 -116.87890625 481.203125 C-114.00360544 480.2446914 -112.58840694 480.13656113 -109.6484375 480.32421875 C-108.84599609 480.37255859 -108.04355469 480.42089844 -107.21679688 480.47070312 C-106.38341797 480.52677734 -105.55003906 480.58285156 -104.69140625 480.640625 C-103.84642578 480.69283203 -103.00144531 480.74503906 -102.13085938 480.79882812 C-100.04654326 480.92836189 -97.96267443 481.06505677 -95.87890625 481.203125 C-98.82308521 478.77983924 -101.96486314 477.06620427 -105.36035156 475.34985352 C-120.5953521 467.64385837 -134.65699067 457.98212651 -147.87890625 447.203125 C-148.4296582 446.75533691 -148.98041016 446.30754883 -149.54785156 445.84619141 C-162.91384059 434.89064997 -175.30255235 422.89713546 -185.87890625 409.203125 C-187.0390625 407.76839844 -187.0390625 407.76839844 -188.22265625 406.3046875 C-214.65281561 373.09970881 -231.30026865 333.27902605 -238.06640625 291.515625 C-238.23325928 290.49525146 -238.4001123 289.47487793 -238.57202148 288.42358398 C-240.5251156 275.90068593 -241.11601326 263.43033484 -241.12890625 250.765625 C-241.12991333 250.06924927 -241.13092041 249.37287354 -241.13195801 248.65539551 C-241.11996634 236.29621671 -240.09260759 224.3665551 -237.87890625 212.203125 C-237.7396875 211.38021973 -237.60046875 210.55731445 -237.45703125 209.70947266 C-230.32233539 167.65275276 -211.75006347 126.63892261 -183.87890625 94.203125 C-183.00413545 93.14672084 -182.13052868 92.08935216 -181.2578125 91.03125 C-170.61476341 78.24084 -159.07005693 66.38078005 -145.87890625 56.203125 C-144.89921875 55.41808594 -143.91953125 54.63304687 -142.91015625 53.82421875 C-116.67404765 32.94476898 -85.58064773 16.58405429 -53.06640625 8.203125 C-52.08591309 7.94893799 -51.10541992 7.69475098 -50.09521484 7.43286133 C-33.66600895 3.278968 -16.98060241 0.08662358 0 0 Z " fill="#F2F1F1" transform="translate(495.87890625,224.796875)"/>
<path d="M0 0 C0.92141785 -0.00701431 1.84283569 -0.01402863 2.79217529 -0.02125549 C5.75603156 -0.03869159 8.71968804 -0.04510954 11.68359375 -0.046875 C13.20199356 -0.04788712 13.20199356 -0.04788712 14.75106812 -0.04891968 C29.7752844 -0.03298984 44.31596387 0.44362914 59.12109375 3.203125 C60.08063965 3.36941406 61.04018555 3.53570312 62.02880859 3.70703125 C84.02343127 7.56010384 105.06616841 14.38909993 125.12109375 24.203125 C126.01151367 24.63608887 126.90193359 25.06905273 127.81933594 25.51513672 C186.52710837 54.34717607 235.36620413 106.64948816 257.05859375 168.765625 C258.11740692 171.90010402 259.13367147 175.04548209 260.12109375 178.203125 C260.32814941 178.86135254 260.53520508 179.51958008 260.74853516 180.19775391 C264.32069212 191.714725 266.70564405 203.45778078 268.74609375 215.328125 C268.86927979 216.03163086 268.99246582 216.73513672 269.11938477 217.45996094 C275.30584129 254.68985964 271.29642037 296.86104155 258.12109375 332.203125 C257.79157715 333.09854004 257.46206055 333.99395508 257.12255859 334.91650391 C248.96730591 356.8174475 239.02469021 377.37167156 225.12109375 396.203125 C224.33001305 397.30026525 223.53962365 398.39790438 222.75 399.49609375 C217.91405607 406.10884897 212.67752814 412.19172125 207.12109375 418.203125 C205.66179636 419.8481036 204.20347065 421.49394469 202.74609375 423.140625 C194.49206878 432.28310405 185.85157861 440.64607322 176.12109375 448.203125 C175.5585791 448.64736816 174.99606445 449.09161133 174.41650391 449.54931641 C145.97735913 471.94869685 113.26113681 488.11313987 78.18676758 497.17700195 C75.58718686 497.85019672 75.58718686 497.85019672 72.12109375 499.203125 C70.97422075 501.2000588 70.97422075 501.2000588 70.12109375 503.203125 C65.92963909 505.13300341 60.59575896 504.24734434 56.05273438 504.1640625 C52.16043789 504.12028784 48.98676122 504.42999151 45.12109375 505.203125 C44.79109375 514.443125 44.46109375 523.683125 44.12109375 533.203125 C45.11109375 533.533125 46.10109375 533.863125 47.12109375 534.203125 C46.46109375 534.533125 45.80109375 534.863125 45.12109375 535.203125 C44.79109375 552.033125 44.46109375 568.863125 44.12109375 586.203125 C26.63109375 586.533125 9.14109375 586.863125 -8.87890625 587.203125 C-9.20890625 604.363125 -9.53890625 621.523125 -9.87890625 639.203125 C-45.18890625 639.203125 -80.49890625 639.203125 -116.87890625 639.203125 C-116.87890625 622.043125 -116.87890625 604.883125 -116.87890625 587.203125 C-134.69890625 586.873125 -152.51890625 586.543125 -170.87890625 586.203125 C-170.89953125 577.64375 -170.92015625 569.084375 -170.94140625 560.265625 C-170.95051025 557.55996338 -170.95961426 554.85430176 -170.96899414 552.06665039 C-170.9719131 549.93636118 -170.9744617 547.80607142 -170.9765625 545.67578125 C-170.98167847 544.55812378 -170.98679443 543.44046631 -170.99206543 542.28894043 C-170.9922467 540.70550842 -170.9922467 540.70550842 -170.99243164 539.09008789 C-170.99465225 538.16853409 -170.99687286 537.24698029 -170.99916077 536.29750061 C-170.87890625 534.203125 -170.87890625 534.203125 -169.87890625 533.203125 C-168.22152182 533.10965585 -166.56015981 533.08567523 -164.90014648 533.08959961 C-163.83912216 533.08967514 -162.77809784 533.08975067 -161.68492126 533.08982849 C-160.53077225 533.09498978 -159.37662323 533.10015106 -158.1875 533.10546875 C-157.01252457 533.1068837 -155.83754913 533.10829865 -154.62696838 533.10975647 C-150.85675561 533.11537508 -147.08660121 533.12793074 -143.31640625 533.140625 C-140.76757898 533.1456376 -138.21875078 533.15020092 -135.66992188 533.15429688 C-129.40620916 533.16450169 -123.14262341 533.18407348 -116.87890625 533.203125 C-116.87890625 516.043125 -116.87890625 498.883125 -116.87890625 481.203125 C-114.00360544 480.2446914 -112.58840694 480.13656113 -109.6484375 480.32421875 C-108.84599609 480.37255859 -108.04355469 480.42089844 -107.21679688 480.47070312 C-106.38341797 480.52677734 -105.55003906 480.58285156 -104.69140625 480.640625 C-103.84642578 480.69283203 -103.00144531 480.74503906 -102.13085938 480.79882812 C-100.04654326 480.92836189 -97.96267443 481.06505677 -95.87890625 481.203125 C-98.82308521 478.77983924 -101.96486314 477.06620427 -105.36035156 475.34985352 C-120.5953521 467.64385837 -134.65699067 457.98212651 -147.87890625 447.203125 C-148.4296582 446.75533691 -148.98041016 446.30754883 -149.54785156 445.84619141 C-162.91384059 434.89064997 -175.30255235 422.89713546 -185.87890625 409.203125 C-187.0390625 407.76839844 -187.0390625 407.76839844 -188.22265625 406.3046875 C-214.65281561 373.09970881 -231.30026865 333.27902605 -238.06640625 291.515625 C-238.23325928 290.49525146 -238.4001123 289.47487793 -238.57202148 288.42358398 C-240.5251156 275.90068593 -241.11601326 263.43033484 -241.12890625 250.765625 C-241.12991333 250.06924927 -241.13092041 249.37287354 -241.13195801 248.65539551 C-241.11996634 236.29621671 -240.09260759 224.3665551 -237.87890625 212.203125 C-237.7396875 211.38021973 -237.60046875 210.55731445 -237.45703125 209.70947266 C-230.32233539 167.65275276 -211.75006347 126.63892261 -183.87890625 94.203125 C-183.00413545 93.14672084 -182.13052868 92.08935216 -181.2578125 91.03125 C-170.61476341 78.24084 -159.07005693 66.38078005 -145.87890625 56.203125 C-144.89921875 55.41808594 -143.91953125 54.63304687 -142.91015625 53.82421875 C-116.67404765 32.94476898 -85.58064773 16.58405429 -53.06640625 8.203125 C-52.08591309 7.94893799 -51.10541992 7.69475098 -50.09521484 7.43286133 C-33.66600895 3.278968 -16.98060241 0.08662358 0 0 Z M-87.87890625 32.203125 C-88.59916992 32.5419873 -89.31943359 32.88084961 -90.06152344 33.22998047 C-124.20445281 49.32727966 -156.09135374 73.99575506 -178.58886719 104.46435547 C-179.89736252 106.22800115 -181.23305076 107.96814091 -182.57421875 109.70703125 C-199.04420168 131.29375941 -211.30332047 155.48240682 -219.87890625 181.203125 C-220.2553125 182.33105469 -220.63171875 183.45898438 -221.01953125 184.62109375 C-226.4402957 202.28160014 -229.96150129 220.96510408 -230.1171875 239.44921875 C-230.12693604 240.40987747 -230.13668457 241.37053619 -230.14672852 242.36030579 C-230.39447879 272.48797364 -230.39447879 272.48797364 -225.87890625 302.203125 C-225.57412354 303.52981201 -225.57412354 303.52981201 -225.26318359 304.88330078 C-224.12315026 309.71078313 -222.85258666 314.48493315 -221.45068359 319.24267578 C-220.94682872 320.97023969 -220.48202696 322.7090916 -220.0234375 324.44921875 C-212.10029768 353.05435734 -196.03025924 379.04512398 -177.87890625 402.203125 C-177.44384766 402.75822754 -177.00878906 403.31333008 -176.56054688 403.88525391 C-164.51746016 419.06047673 -150.53862363 432.80514308 -134.87890625 444.203125 C-133.72895794 445.05961566 -132.57922036 445.91638933 -131.4296875 446.7734375 C-118.38213271 456.39532293 -104.52167673 464.28056306 -89.87890625 471.203125 C-89.25999512 471.49928711 -88.64108398 471.79544922 -88.00341797 472.10058594 C-72.22710666 479.58213563 -55.49532469 485.11639531 -38.50390625 489.078125 C-37.69872559 489.26906738 -36.89354492 489.46000977 -36.06396484 489.65673828 C-20.9766374 492.96186682 -5.70493714 493.55482762 9.68359375 493.453125 C10.55471802 493.44935852 11.42584229 493.44559204 12.32336426 493.44171143 C82.57194596 493.08730937 143.90360263 468.03485208 193.50439453 418.05395508 C198.74019809 412.69604669 203.54923926 407.14018604 208.12109375 401.203125 C209.09871795 399.9987463 210.07800766 398.79571841 211.05859375 397.59375 C226.80105761 378.01476626 239.94241947 355.03391103 247.26953125 330.90625 C247.9368453 328.78798706 248.71580523 326.70484636 249.53515625 324.640625 C251.59016263 319.21071973 252.8294667 313.60399336 254.12109375 307.953125 C254.36859375 306.91671875 254.61609375 305.8803125 254.87109375 304.8125 C258.86323226 287.51323312 260.65397018 270.68692135 260.49609375 252.953125 C260.49144104 252.01568451 260.48678833 251.07824402 260.48199463 250.11239624 C260.0975485 183.86162534 232.6354719 125.13103863 185.9230957 78.77075195 C180.58381826 73.55485172 175.06358531 68.72615501 169.12109375 64.203125 C168.5286084 63.74486328 167.93612305 63.28660156 167.32568359 62.81445312 C135.66256562 38.33700882 100.42530512 22.10062248 61.18359375 14.078125 C60.42264404 13.91965088 59.66169434 13.76117676 58.87768555 13.59790039 C44.20000168 10.68863104 29.79537058 9.79010718 14.87109375 9.828125 C13.49114227 9.83043625 13.49114227 9.83043625 12.08331299 9.83279419 C-22.78749818 9.97113752 -56.37350221 17.02799914 -87.87890625 32.203125 Z " fill="#ECECEC" transform="translate(495.87890625,224.796875)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C56.25055952 6.50111903 56.15703468 18.1037619 53.9375 24.97265625 C53.21240669 26.8704897 52.41986391 28.72829718 51.61376953 30.59301758 C44.98617599 46.02400619 42.04821032 63.39466522 40 80 C39.90501221 80.73130127 39.81002441 81.46260254 39.7121582 82.21606445 C38.81242058 89.94101176 38.80128667 97.6689295 38.8125 105.4375 C38.81277191 106.14587006 38.81304382 106.85424011 38.81332397 107.58407593 C38.83315593 118.83799648 39.36546858 129.85844861 41 141 C41.10183594 141.7542627 41.20367187 142.50852539 41.30859375 143.28564453 C42.06463387 148.88477498 42.96797621 154.44518506 44 160 C44.14743652 160.79535156 44.29487305 161.59070313 44.44677734 162.41015625 C51.82214009 200.50218517 70.60781395 236.09841748 95 266 C95.45310547 266.55606934 95.90621094 267.11213867 96.37304688 267.68505859 C107.05024901 280.68004843 118.63626677 292.74329061 132 303 C132.58475098 303.45584473 133.16950195 303.91168945 133.77197266 304.38134766 C143.4650023 311.92644768 153.47406951 318.67324391 164 325 C162.515 330.445 162.515 330.445 161 336 C156.50610584 336.17159991 152.01196957 336.33158549 147.51733398 336.48217773 C145.99802334 336.53455678 144.47880665 336.58976042 142.9597168 336.64819336 C131.18422369 337.09823713 119.83438086 336.62286215 108 336 C107.01 310.26 107.01 310.26 106 284 C88.84 284 71.68 284 54 284 C54 300.83 54 317.66 54 335 C49.71069382 336.71572247 48.21089419 337.24575954 43.93432617 337.13525391 C42.94009644 337.11470947 41.9458667 337.09416504 40.92150879 337.07299805 C39.88909058 337.04117432 38.85667236 337.00935059 37.79296875 336.9765625 C36.35564392 336.94405396 36.35564392 336.94405396 34.88928223 336.91088867 C31.32173236 336.82711225 27.7546329 336.72496711 24.1875 336.625 C16.205625 336.41875 8.22375 336.2125 0 336 C0 318.84 0 301.68 0 284 C-17.82 284 -35.64 284 -54 284 C-55.24177521 281.51644959 -55.12036681 279.86892378 -55.11352539 277.09130859 C-55.11340454 276.05611084 -55.11328369 275.02091309 -55.11315918 273.9543457 C-55.10804321 272.863396 -55.10292725 271.77244629 -55.09765625 270.6484375 C-55.09664917 269.6478833 -55.09564209 268.6473291 -55.09460449 267.61645508 C-55.08936192 263.86929177 -55.07540072 260.12214477 -55.0625 256.375 C-55.041875 248.00125 -55.02125 239.6275 -55 231 C-72.49 231 -89.98 231 -108 231 C-108.020625 222.440625 -108.04125 213.88125 -108.0625 205.0625 C-108.071604 202.35683838 -108.08070801 199.65117676 -108.09008789 196.86352539 C-108.09300685 194.73323618 -108.09555545 192.60294642 -108.09765625 190.47265625 C-108.10277222 189.35499878 -108.10788818 188.23734131 -108.11315918 187.08581543 C-108.11328003 186.03019409 -108.11340088 184.97457275 -108.11352539 183.88696289 C-108.115746 182.96540909 -108.11796661 182.04385529 -108.12025452 181.09437561 C-108 179 -108 179 -107 178 C-105.37325222 177.90659566 -103.74245949 177.88254829 -102.11303711 177.88647461 C-100.5296051 177.88665588 -100.5296051 177.88665588 -98.91418457 177.88684082 C-97.7965271 177.89195679 -96.67886963 177.89707275 -95.52734375 177.90234375 C-93.99551453 177.90385437 -93.99551453 177.90385437 -92.43273926 177.90539551 C-88.60098149 177.91064585 -84.76923967 177.92460697 -80.9375 177.9375 C-72.378125 177.958125 -63.81875 177.97875 -55 178 C-55 160.84 -55 143.68 -55 126 C-61.6 126 -68.2 126 -75 126 C-80.91869453 125.85883863 -86.83352956 125.70094691 -92.75 125.5 C-94.24868845 125.45152929 -95.74738641 125.40335181 -97.24609375 125.35546875 C-100.83084412 125.24032449 -104.41545315 125.12133504 -108 125 C-108.02888146 121.68751813 -108.04675799 118.37506833 -108.0625 115.0625 C-108.07087891 114.11697266 -108.07925781 113.17144531 -108.08789062 112.19726562 C-108.09111328 111.29814453 -108.09433594 110.39902344 -108.09765625 109.47265625 C-108.10289307 108.64000244 -108.10812988 107.80734863 -108.11352539 106.94946289 C-108 105 -108 105 -107 104 C-105.41484422 103.89625042 -103.82510534 103.86148111 -102.23657227 103.85473633 C-101.22204483 103.84835648 -100.2075174 103.84197662 -99.1622467 103.83540344 C-98.05811935 103.83429062 -96.953992 103.8331778 -95.81640625 103.83203125 C-94.12764626 103.82703865 -94.12764626 103.82703865 -92.4047699 103.82194519 C-90.01814179 103.81687106 -87.63150655 103.81453701 -85.24487305 103.81469727 C-81.58175026 103.81251149 -77.91892878 103.7943626 -74.25585938 103.77539062 C-71.94270937 103.77245674 -69.62955792 103.77047191 -67.31640625 103.76953125 C-66.21430313 103.76234573 -65.11220001 103.75516022 -63.97669983 103.74775696 C-62.45018044 103.7523719 -62.45018044 103.7523719 -60.89282227 103.75708008 C-59.99427017 103.75565506 -59.09571808 103.75423004 -58.16993713 103.75276184 C-56 104 -56 104 -54 106 C-54 112.6 -54 119.2 -54 126 C-35.85 126 -17.7 126 1 126 C0.67 125.67 0.34 125.34 0 125 C-0.495 114.605 -0.495 114.605 -1 104 C-18.49 104 -35.98 104 -54 104 C-54 87.17 -54 70.34 -54 53 C-46.48856893 52.97708377 -38.97725844 52.95715862 -31.46582031 52.94506836 C-28.90884999 52.94002983 -26.35188257 52.93319893 -23.79492188 52.92456055 C-20.12629483 52.91247398 -16.45770577 52.90676699 -12.7890625 52.90234375 C-11.64007477 52.89718246 -10.49108704 52.89202118 -9.30728149 52.88670349 C-8.2463327 52.88662796 -7.18538391 52.88655243 -6.09228516 52.88647461 C-5.15518707 52.884254 -4.21808899 52.88203339 -3.25259399 52.87974548 C-1 53 -1 53 1 54 C0.67 53.34 0.34 52.68 0 52 C-0.09039906 50.3351936 -0.11755257 48.66676579 -0.11352539 46.99951172 C-0.11340454 45.94401123 -0.11328369 44.88851074 -0.11315918 43.80102539 C-0.10804321 42.68848389 -0.10292725 41.57594238 -0.09765625 40.4296875 C-0.09664917 39.4094751 -0.09564209 38.3892627 -0.09460449 37.33813477 C-0.08936163 33.51707845 -0.07540043 29.69603813 -0.0625 25.875 C-0.041875 17.33625 -0.02125 8.7975 0 0 Z " fill="#F8F8F8" transform="translate(217,369)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C3.31303391 13.57754211 -0.52046332 25.68900446 -4.5 37.5 C-4.71586761 38.14241638 -4.93173523 38.78483276 -5.15414429 39.44671631 C-15.72995012 70.70214139 -32.78378295 97.72481583 -55.55322266 121.48583984 C-56.91633676 122.9124402 -58.26153241 124.35610006 -59.60546875 125.80078125 C-67.32056227 133.8660303 -75.9754894 140.47180916 -85 147 C-85.61327148 147.44730469 -86.22654297 147.89460937 -86.85839844 148.35546875 C-102.91896159 159.94832389 -120.86037412 169.01284916 -139.65454102 175.21777344 C-141.34975554 175.78313904 -143.0369131 176.37286035 -144.71850586 176.97753906 C-152.43954969 179.69862306 -160.12753972 181.3668012 -168.1875 182.75 C-169.99637695 183.08064453 -169.99637695 183.08064453 -171.84179688 183.41796875 C-178.32976745 184.55894446 -184.41411861 185.25466351 -191 185 C-190.98428955 185.59014893 -190.9685791 186.18029785 -190.95239258 186.78833008 C-190.89002061 189.46295586 -190.85100343 192.13742864 -190.8125 194.8125 C-190.78736328 195.74126953 -190.76222656 196.67003906 -190.73632812 197.62695312 C-190.72666016 198.51962891 -190.71699219 199.41230469 -190.70703125 200.33203125 C-190.6913208 201.15421143 -190.67561035 201.9763916 -190.65942383 202.82348633 C-191.08015812 205.512265 -191.83123218 206.39977562 -194 208 C-197.22319552 207.9217671 -198.70080292 207.24157785 -201.2109375 205.21484375 C-201.92507813 204.46332031 -202.63921875 203.71179688 -203.375 202.9375 C-204.08398438 202.20402344 -204.79296875 201.47054687 -205.5234375 200.71484375 C-207.42236809 198.63320849 -209.26360713 196.52785386 -211.09692383 194.38989258 C-215.17002099 189.73083795 -219.5197858 185.38899588 -223.92578125 181.046875 C-225.62578147 179.35950639 -227.32564739 177.67200248 -229.02539062 175.984375 C-231.68113538 173.35354713 -234.33846515 170.7243582 -236.99829102 168.09765625 C-239.58265063 165.5434218 -242.16081925 162.98306692 -244.73828125 160.421875 C-245.53720291 159.63641296 -246.33612457 158.85095093 -247.15925598 158.04168701 C-247.89729965 157.30702209 -248.63534332 156.57235718 -249.39575195 155.81542969 C-250.04526321 155.17337585 -250.69477448 154.53132202 -251.3639679 153.86981201 C-255.05847966 149.64737503 -255.77401315 145.57705502 -255.59747314 140.0632019 C-254.87701811 136.36948068 -253.70523891 135.00476647 -251.11621094 132.30908203 C-250.2965686 131.4449469 -249.47692627 130.58081177 -248.63244629 129.69049072 C-247.76373901 128.80262878 -246.89503174 127.91476685 -246 127 C-245.17028687 126.13614685 -244.34057373 125.2722937 -243.48571777 124.38226318 C-237.83868821 118.53791219 -232.09961353 112.78247034 -226.36962891 107.01953125 C-224.27566865 104.91210448 -222.18927548 102.79758173 -220.10888672 100.67675781 C-217.57433788 98.09300089 -215.02783217 95.52163489 -212.47212982 92.95880508 C-211.50622674 91.98619557 -210.54457832 91.00934094 -209.58737946 90.02816391 C-208.25527773 88.66453408 -206.9058279 87.31791644 -205.55566406 85.97216797 C-204.7944928 85.20290985 -204.03332153 84.43365173 -203.24908447 83.64108276 C-200.57116415 81.68709262 -199.24412347 81.55345952 -196 82 C-194.20581055 83.15356445 -194.20581055 83.15356445 -193 85 C-192.65942383 87.54370117 -192.65942383 87.54370117 -192.70703125 90.54296875 C-192.7215332 92.15268555 -192.7215332 92.15268555 -192.73632812 93.79492188 C-192.76146484 94.91447266 -192.78660156 96.03402344 -192.8125 97.1875 C-192.83280273 98.88422852 -192.83280273 98.88422852 -192.85351562 100.61523438 C-192.88890042 103.41063317 -192.93827052 106.20507892 -193 109 C-156.53250316 101.25829676 -122.75293558 81.97157126 -101.65234375 50.59375 C-96.40003038 42.34898386 -91.84149486 33.99299257 -88 25 C-85.14447237 26.2979671 -83.11891706 27.69873873 -80.875 29.875 C-72.47036503 37.31546689 -61.78707553 38.65488546 -51 38 C-39.10718265 36.11855284 -30.0801439 28.43126638 -21.56640625 20.4140625 C-19.34572474 18.32520227 -17.07896896 16.34048826 -14.75 14.375 C-11.27073159 11.37538382 -8.34652287 8.0595757 -5.4453125 4.50390625 C-4.96835937 4.00761719 -4.49140625 3.51132812 -4 3 C-3.34 3 -2.68 3 -2 3 C-2 2.34 -2 1.68 -2 1 C-1.34 0.67 -0.68 0.34 0 0 Z " fill="#E26A98" transform="translate(729,498)"/>
<path d="M0 0 C13.91724179 -1.78087928 13.91724179 -1.78087928 18.98291016 1.14550781 C22.89053317 4.27538475 26.08493024 7.94473917 29 12 C29 12.66 29 13.32 29 14 C29.66 14 30.32 14 31 14 C32.27172852 15.3215332 32.27172852 15.3215332 33.81640625 17.23828125 C37.04016932 21.04043272 40.49972899 24.41627848 44.15234375 27.79296875 C45.84013186 29.38322658 47.52482236 30.97671773 49.20922852 32.57055664 C50.36367905 33.65064223 51.52853939 34.71970511 52.70336914 35.77758789 C63.72764161 45.74475939 63.72764161 45.74475939 64.19140625 53.80078125 C64.01221476 60.27309436 60.29077623 63.59701311 56 68 C55.2638295 68.76147842 54.527659 69.52295685 53.7691803 70.30751038 C51.27567088 72.85643005 48.75866123 75.38000328 46.234375 77.8984375 C45.31916077 78.81460846 44.40394653 79.73077942 43.46099854 80.67471313 C41.53974333 82.5974303 39.61672231 84.51835817 37.69238281 86.43798828 C35.22880501 88.89582921 32.76979914 91.35818799 30.31206894 93.82187462 C27.9552631 96.18315876 25.5946596 98.5406306 23.234375 100.8984375 C22.35311951 101.78171722 21.47186401 102.66499695 20.56390381 103.57504272 C19.74585266 104.38994171 18.92780151 105.2048407 18.08496094 106.04443359 C17.36661072 106.76198822 16.6482605 107.47954285 15.90814209 108.21884155 C13.00920304 110.92486109 11.44897267 111.96061643 7.4375 112.3125 C6.303125 112.209375 5.16875 112.10625 4 112 C1.76586987 108.64880481 1.76152238 107.5822245 1.8046875 103.67578125 C1.81435547 102.13374023 1.81435547 102.13374023 1.82421875 100.56054688 C1.84935547 98.95276367 1.84935547 98.95276367 1.875 97.3125 C1.88402344 96.22904297 1.89304687 95.14558594 1.90234375 94.02929688 C1.9259266 91.3526429 1.95883874 88.67643203 2 86 C-33.60229911 93.005082 -65.00644976 110.71227547 -86 141 C-92.60895162 150.89119005 -98.40061183 161.01580716 -103 172 C-103.94875 171.13375 -104.8975 170.2675 -105.875 169.375 C-115.5010328 161.15195174 -124.65395632 157.39964714 -137.37109375 157.62890625 C-152.26554967 159.15202069 -162.25433757 170.0591707 -172.17578125 180.171875 C-175.06909724 183.06919281 -178.06370957 185.75623143 -181.1875 188.3984375 C-183.77298557 190.68302604 -186.11498117 193.18364948 -188.45703125 195.71484375 C-190 197 -190 197 -193 197 C-193.16898963 190.69731283 -192.68400316 185.08124149 -191.3125 178.9375 C-191.13388428 178.11822021 -190.95526855 177.29894043 -190.77124023 176.45483398 C-186.66718315 158.21320853 -179.61826837 141.5321212 -171 125 C-170.66516602 124.35015137 -170.33033203 123.70030273 -169.98535156 123.03076172 C-161.77745158 107.23869859 -151.21408254 92.923919 -139 80 C-137.78572343 78.60933378 -136.57714048 77.21367037 -135.375 75.8125 C-128.86482247 68.38079049 -121.73856811 62.14060404 -114 56 C-112.98679687 55.18144531 -111.97359375 54.36289062 -110.9296875 53.51953125 C-103.04356367 47.22603286 -94.77008971 41.97017286 -86 37 C-85.41025391 36.65727051 -84.82050781 36.31454102 -84.21289062 35.96142578 C-59.65651517 21.72772203 -28.54389817 11.14794334 0 12 C0 8.04 0 4.08 0 0 Z " fill="#2ECC9C" transform="translate(484,259)"/>
<path d="M0 0 C7.40084051 -0.45348287 13.87847358 1.21315092 21 3.125 C22.20897949 3.44702393 23.41795898 3.76904785 24.66357422 4.10083008 C47.73887755 10.36863575 70.4435235 20.10186404 90 34 C91.45019531 35.01513672 91.45019531 35.01513672 92.9296875 36.05078125 C138.99748006 68.91077179 170.22887434 115.65403091 180.73828125 171.3828125 C181.12540351 175.25403513 181.05227103 179.11293647 181 183 C181.62567871 182.98952637 182.25135742 182.97905273 182.89599609 182.96826172 C185.7222901 182.92676809 188.54852011 182.90069527 191.375 182.875 C192.35984375 182.85824219 193.3446875 182.84148437 194.359375 182.82421875 C195.30039062 182.81777344 196.24140625 182.81132812 197.2109375 182.8046875 C198.51490479 182.78897705 198.51490479 182.78897705 199.84521484 182.77294922 C202 183 202 183 204 185 C204.5 187.1875 204.5 187.1875 204 190 C202.25247516 192.58376373 200.32164007 194.91292979 198 197 C197.34 197 196.68 197 196 197 C196 197.66 196 198.32 196 199 C194.51367188 200.46508789 194.51367188 200.46508789 192.46875 202.16015625 C188.26922235 205.73326051 184.37163803 209.51515257 180.5 213.4375 C179.82001953 214.12126709 179.14003906 214.80503418 178.43945312 215.50952148 C176.29049074 217.67057055 174.14482721 219.83484726 172 222 C169.16966163 224.85716017 166.33587327 227.71083454 163.5 230.5625 C162.54963867 231.52530884 162.54963867 231.52530884 161.58007812 232.50756836 C145.76825224 248.40442636 145.76825224 248.40442636 138.75 248.625 C137.85796875 248.67914063 136.9659375 248.73328125 136.046875 248.7890625 C124.20354617 245.72194401 112.18257248 228.52645634 103.46142578 219.86645508 C101.14747312 217.57042989 98.82526297 215.2832607 96.49560547 213.00317383 C93.66555142 210.23322412 90.85042392 207.44890924 88.04541016 204.65361214 C86.97878063 203.59553454 85.90702879 202.54259426 84.83007812 201.49502373 C83.32934108 200.03312137 81.84856689 198.55347475 80.37109375 197.06811523 C79.52474365 196.2320726 78.67839355 195.39602997 77.80639648 194.53465271 C75.58912981 191.42348578 75.46921807 189.74331841 76 186 C78 184 78 184 80.43017578 183.77294922 C81.92266846 183.78865967 81.92266846 183.78865967 83.4453125 183.8046875 C85.05986328 183.81435547 85.05986328 183.81435547 86.70703125 183.82421875 C87.83496094 183.84097656 88.96289062 183.85773438 90.125 183.875 C91.26066406 183.88402344 92.39632812 183.89304687 93.56640625 183.90234375 C96.37781299 183.92596902 99.18880298 183.95890987 102 184 C97.58956696 164.17733086 89.71760425 145.93023947 77 130 C76.35853027 129.18233154 76.35853027 129.18233154 75.70410156 128.34814453 C68.42269641 119.1371927 60.55933299 111.79229225 51 105 C50.08879395 104.34257812 50.08879395 104.34257812 49.15917969 103.671875 C40.23968819 97.28403486 31.07771345 92.31697796 21 88 C22.18883856 84.67575948 23.33065668 82.37648852 25.8125 79.875 C33.36061531 71.17704894 34.93571908 62.43455472 34.41015625 51.2421875 C33.98940244 45.89544966 32.77294066 41.61359955 30 37 C29.51015625 36.18144531 29.0203125 35.36289062 28.515625 34.51953125 C23.28401454 26.68368992 16.53434483 20.33168338 9.8046875 13.796875 C2.22837 6.33887783 2.22837 6.33887783 0 3 C0 2.01 0 1.02 0 0 Z " fill="#E54176" transform="translate(539,263)"/>
<path d="M0 0 C1.89355469 1.21704102 1.89355469 1.21704102 3.671875 2.87890625 C4.35668945 3.51449463 5.04150391 4.15008301 5.74707031 4.80493164 C10.97045754 9.89416816 16.10290617 15.06851458 21.22265625 20.26171875 C25.77729857 24.8561396 30.35179293 29.32212291 35.30786133 33.48388672 C37.60594864 35.54291459 39.54545865 37.8297222 41.48046875 40.2265625 C44.32148228 43.54229551 47.46200285 46.51781812 50.7109375 49.4296875 C51.59007812 50.23664063 52.46921875 51.04359375 53.375 51.875 C54.26960938 52.67679687 55.16421875 53.47859375 56.0859375 54.3046875 C58 57 58 57 57.9140625 60.7578125 C57.61242187 61.82773437 57.31078125 62.89765625 57 64 C54.44276771 65.27861615 52.63262898 65.11336609 49.7734375 65.09765625 C48.2265625 65.09282227 48.2265625 65.09282227 46.6484375 65.08789062 C45.56820312 65.07951172 44.48796875 65.07113281 43.375 65.0625 C41.74304688 65.05573242 41.74304688 65.05573242 40.078125 65.04882812 C37.38536211 65.03701776 34.69270812 65.02054778 32 65 C38.32332591 96.73445549 55.61317907 124.36923361 82.38671875 143.07421875 C91.72932816 149.23636538 101.98605359 154.03997646 112 159 C112 163.69475512 111.46939999 163.96226471 108.3125 167.125 C99.91480387 176.14805648 97.5374923 185.18801335 97.6640625 197.30078125 C99.03324574 212.37771759 110.30794023 222.57461124 120.54443359 232.55981445 C129.55989554 241.36925579 129.55989554 241.36925579 132 245 C132 245.99 132 246.98 132 248 C124.80430205 248.40121467 118.50291191 246.95042886 111.5625 245.125 C110.37962402 244.81401367 109.19674805 244.50302734 107.97802734 244.18261719 C82.52531399 237.2258809 58.05893205 226.02362912 36.79833984 210.32666016 C35.64438509 209.47537179 34.48373945 208.63303763 33.31494141 207.80224609 C16.59799833 195.91563807 0.55918977 179.94914904 -11 163 C-11.84100572 161.80328694 -12.6821585 160.60667721 -13.5234375 159.41015625 C-32.23425204 132.42785676 -46.61782282 98.22895229 -46 65 C-46.65597168 65.01047363 -47.31194336 65.02094727 -47.98779297 65.03173828 C-50.95015658 65.07322503 -53.91245916 65.09930262 -56.875 65.125 C-57.90753906 65.14175781 -58.94007813 65.15851563 -60.00390625 65.17578125 C-60.99003906 65.18222656 -61.97617187 65.18867188 -62.9921875 65.1953125 C-63.90339355 65.20578613 -64.81459961 65.21625977 -65.75341797 65.22705078 C-68 65 -68 65 -70 63 C-70.09041316 59.53122833 -69.81579918 57.04576542 -67.63516235 54.25042725 C-65.71312289 52.35001152 -63.72025991 50.5727787 -61.67578125 48.8046875 C-60.11244486 47.39486844 -58.55218686 45.98163012 -56.99462891 44.56542969 C-56.17496643 43.82417847 -55.35530396 43.08292725 -54.51080322 42.31921387 C-50.27109637 38.40302209 -46.22366887 34.30042293 -42.16796875 30.1953125 C-41.34861847 29.36997009 -40.52926819 28.54462769 -39.68508911 27.6942749 C-36.31972541 24.30331516 -32.9596667 20.90716073 -29.60327148 17.50732422 C-27.10832759 14.98232646 -24.60731067 12.46347288 -22.10546875 9.9453125 C-20.96962593 8.78928024 -20.96962593 8.78928024 -19.81083679 7.6098938 C-19.1052211 6.90089935 -18.39960541 6.19190491 -17.67260742 5.46142578 C-17.05769943 4.83906036 -16.44279144 4.21669495 -15.80924988 3.57546997 C-11.04981603 -0.56897973 -6.08106451 -1.05528234 0 0 Z " fill="#804D8B" transform="translate(350,442)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.90744461 0.00680466 4.96846893 0.00688019 6.06164551 0.00695801 C7.21579453 0.01211929 8.36994354 0.01728058 9.55906677 0.02259827 C10.73404221 0.02401321 11.90901764 0.02542816 13.11959839 0.02688599 C16.88981116 0.0325046 20.65996556 0.04506026 24.43016052 0.05775452 C26.97898779 0.06276712 29.52781599 0.06733044 32.0766449 0.07142639 C38.34033685 0.08248007 44.60399452 0.0992363 50.86766052 0.12025452 C51.01282423 5.11488994 51.1550925 10.10959733 51.29490662 15.10438538 C51.34265205 16.7964642 51.39113026 18.48852254 51.44041443 20.18055725 C51.68838271 28.71016003 51.91524212 37.23915994 51.96141052 45.77259827 C51.96850037 46.97779114 51.97559021 48.18298401 51.9828949 49.42469788 C51.86766052 52.12025452 51.86766052 52.12025452 50.86766052 53.12025452 C49.21121686 53.2431617 47.5496706 53.29809359 45.88890076 53.32557678 C44.82787643 53.345522 43.76685211 53.36546722 42.67367554 53.38601685 C41.51952652 53.40272934 40.3653775 53.41944183 39.17625427 53.43666077 C38.00127884 53.45744186 36.82630341 53.47822296 35.61572266 53.49963379 C31.84559729 53.56525576 28.0753997 53.62407282 24.30516052 53.68275452 C21.75632479 53.72592772 19.20749649 53.7695416 16.65867615 53.81361389 C10.39507734 53.92178292 4.13142733 54.02076245 -2.13233948 54.12025452 C-2.46233948 71.28025452 -2.79233948 88.44025452 -3.13233948 106.12025452 C14.68766052 106.12025452 32.50766052 106.12025452 50.86766052 106.12025452 C50.82874165 96.90903966 50.82874165 96.90903966 50.77757263 87.69789124 C50.75353392 76.1112344 51.33934764 64.74313786 51.86766052 53.12025452 C69.35766052 53.12025452 86.84766052 53.12025452 104.86766052 53.12025452 C104.86766052 70.61025452 104.86766052 88.10025452 104.86766052 106.12025452 C87.37766052 106.45025452 69.88766052 106.78025452 51.86766052 107.12025452 C51.53766052 123.95025452 51.20766052 140.78025452 50.86766052 158.12025452 C33.04766052 158.12025452 15.22766052 158.12025452 -3.13233948 158.12025452 C-3.13233948 175.61025452 -3.13233948 193.10025452 -3.13233948 211.12025452 C-20.62233948 211.12025452 -38.11233948 211.12025452 -56.13233948 211.12025452 C-56.13233948 193.63025452 -56.13233948 176.14025452 -56.13233948 158.12025452 C-73.95233948 158.12025452 -91.77233948 158.12025452 -110.13233948 158.12025452 C-110.13233948 140.96025452 -110.13233948 123.80025452 -110.13233948 106.12025452 C-92.31233948 106.12025452 -74.49233948 106.12025452 -56.13233948 106.12025452 C-56.13233948 88.63025452 -56.13233948 71.14025452 -56.13233948 53.12025452 C-38.64233948 53.12025452 -21.15233948 53.12025452 -3.13233948 53.12025452 C-3.17194918 36.05200152 -3.17194918 36.05200152 -3.22242737 18.98377991 C-3.22534633 16.8534907 -3.22789493 14.72320094 -3.22999573 12.59291077 C-3.23511169 11.4752533 -3.24022766 10.35759583 -3.24549866 9.20606995 C-3.24567993 7.62263794 -3.24567993 7.62263794 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#EFEFEF" transform="translate(758.1323394775391,52.87974548339844)"/>
<path d="M0 0 C0.92141785 -0.00701431 1.84283569 -0.01402863 2.79217529 -0.02125549 C5.75603156 -0.03869159 8.71968804 -0.04510954 11.68359375 -0.046875 C13.20199356 -0.04788712 13.20199356 -0.04788712 14.75106812 -0.04891968 C29.7752844 -0.03298984 44.31596387 0.44362914 59.12109375 3.203125 C60.08063965 3.36941406 61.04018555 3.53570312 62.02880859 3.70703125 C84.02343127 7.56010384 105.06616841 14.38909993 125.12109375 24.203125 C126.01151367 24.63608887 126.90193359 25.06905273 127.81933594 25.51513672 C186.52710837 54.34717607 235.36620413 106.64948816 257.05859375 168.765625 C258.11740692 171.90010402 259.13367147 175.04548209 260.12109375 178.203125 C260.32814941 178.86135254 260.53520508 179.51958008 260.74853516 180.19775391 C264.32069212 191.714725 266.70564405 203.45778078 268.74609375 215.328125 C268.86927979 216.03163086 268.99246582 216.73513672 269.11938477 217.45996094 C275.30584129 254.68985964 271.29642037 296.86104155 258.12109375 332.203125 C257.79157715 333.09854004 257.46206055 333.99395508 257.12255859 334.91650391 C248.96730591 356.8174475 239.02469021 377.37167156 225.12109375 396.203125 C224.33001305 397.30026525 223.53962365 398.39790438 222.75 399.49609375 C217.91405607 406.10884897 212.67752814 412.19172125 207.12109375 418.203125 C205.66179636 419.8481036 204.20347065 421.49394469 202.74609375 423.140625 C194.49206878 432.28310405 185.85157861 440.64607322 176.12109375 448.203125 C175.5585791 448.64736816 174.99606445 449.09161133 174.41650391 449.54931641 C138.82208495 477.58436944 96.85970836 495.44446233 52.12109375 502.203125 C50.93531738 502.38319092 50.93531738 502.38319092 49.72558594 502.56689453 C-17.4429433 512.1359143 -85.85804337 493.90239448 -140.03662109 453.41748047 C-142.68977026 451.3940576 -145.29301086 449.31124391 -147.87890625 447.203125 C-148.4296582 446.75533691 -148.98041016 446.30754883 -149.54785156 445.84619141 C-162.91384059 434.89064997 -175.30255235 422.89713546 -185.87890625 409.203125 C-187.0390625 407.76839844 -187.0390625 407.76839844 -188.22265625 406.3046875 C-214.65281561 373.09970881 -231.30026865 333.27902605 -238.06640625 291.515625 C-238.23325928 290.49525146 -238.4001123 289.47487793 -238.57202148 288.42358398 C-240.5251156 275.90068593 -241.11601326 263.43033484 -241.12890625 250.765625 C-241.12991333 250.06924927 -241.13092041 249.37287354 -241.13195801 248.65539551 C-241.11996634 236.29621671 -240.09260759 224.3665551 -237.87890625 212.203125 C-237.7396875 211.38021973 -237.60046875 210.55731445 -237.45703125 209.70947266 C-230.32233539 167.65275276 -211.75006347 126.63892261 -183.87890625 94.203125 C-183.00413545 93.14672084 -182.13052868 92.08935216 -181.2578125 91.03125 C-170.61476341 78.24084 -159.07005693 66.38078005 -145.87890625 56.203125 C-144.89921875 55.41808594 -143.91953125 54.63304687 -142.91015625 53.82421875 C-116.67404765 32.94476898 -85.58064773 16.58405429 -53.06640625 8.203125 C-52.08591309 7.94893799 -51.10541992 7.69475098 -50.09521484 7.43286133 C-33.66600895 3.278968 -16.98060241 0.08662358 0 0 Z M-87.87890625 32.203125 C-88.59916992 32.5419873 -89.31943359 32.88084961 -90.06152344 33.22998047 C-124.20445281 49.32727966 -156.09135374 73.99575506 -178.58886719 104.46435547 C-179.89736252 106.22800115 -181.23305076 107.96814091 -182.57421875 109.70703125 C-199.04420168 131.29375941 -211.30332047 155.48240682 -219.87890625 181.203125 C-220.2553125 182.33105469 -220.63171875 183.45898438 -221.01953125 184.62109375 C-226.4402957 202.28160014 -229.96150129 220.96510408 -230.1171875 239.44921875 C-230.12693604 240.40987747 -230.13668457 241.37053619 -230.14672852 242.36030579 C-230.39447879 272.48797364 -230.39447879 272.48797364 -225.87890625 302.203125 C-225.57412354 303.52981201 -225.57412354 303.52981201 -225.26318359 304.88330078 C-224.12315026 309.71078313 -222.85258666 314.48493315 -221.45068359 319.24267578 C-220.94682872 320.97023969 -220.48202696 322.7090916 -220.0234375 324.44921875 C-212.10029768 353.05435734 -196.03025924 379.04512398 -177.87890625 402.203125 C-177.44384766 402.75822754 -177.00878906 403.31333008 -176.56054688 403.88525391 C-164.51746016 419.06047673 -150.53862363 432.80514308 -134.87890625 444.203125 C-133.72895794 445.05961566 -132.57922036 445.91638933 -131.4296875 446.7734375 C-118.38213271 456.39532293 -104.52167673 464.28056306 -89.87890625 471.203125 C-89.25999512 471.49928711 -88.64108398 471.79544922 -88.00341797 472.10058594 C-72.22710666 479.58213563 -55.49532469 485.11639531 -38.50390625 489.078125 C-37.69872559 489.26906738 -36.89354492 489.46000977 -36.06396484 489.65673828 C-20.9766374 492.96186682 -5.70493714 493.55482762 9.68359375 493.453125 C10.55471802 493.44935852 11.42584229 493.44559204 12.32336426 493.44171143 C82.57194596 493.08730937 143.90360263 468.03485208 193.50439453 418.05395508 C198.74019809 412.69604669 203.54923926 407.14018604 208.12109375 401.203125 C209.09871795 399.9987463 210.07800766 398.79571841 211.05859375 397.59375 C226.80105761 378.01476626 239.94241947 355.03391103 247.26953125 330.90625 C247.9368453 328.78798706 248.71580523 326.70484636 249.53515625 324.640625 C251.59016263 319.21071973 252.8294667 313.60399336 254.12109375 307.953125 C254.36859375 306.91671875 254.61609375 305.8803125 254.87109375 304.8125 C258.86323226 287.51323312 260.65397018 270.68692135 260.49609375 252.953125 C260.49144104 252.01568451 260.48678833 251.07824402 260.48199463 250.11239624 C260.0975485 183.86162534 232.6354719 125.13103863 185.9230957 78.77075195 C180.58381826 73.55485172 175.06358531 68.72615501 169.12109375 64.203125 C168.5286084 63.74486328 167.93612305 63.28660156 167.32568359 62.81445312 C135.66256562 38.33700882 100.42530512 22.10062248 61.18359375 14.078125 C60.42264404 13.91965088 59.66169434 13.76117676 58.87768555 13.59790039 C44.20000168 10.68863104 29.79537058 9.79010718 14.87109375 9.828125 C13.49114227 9.83043625 13.49114227 9.83043625 12.08331299 9.83279419 C-22.78749818 9.97113752 -56.37350221 17.02799914 -87.87890625 32.203125 Z " fill="#16504E" transform="translate(495.87890625,224.796875)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C71.06825299 51.9603903 71.06825299 51.9603903 88.13647461 51.90991211 C90.26676382 51.90699315 92.39705358 51.90444455 94.52734375 51.90234375 C95.64500122 51.89722778 96.76265869 51.89211182 97.91418457 51.88684082 C99.49761658 51.88665955 99.49761658 51.88665955 101.11303711 51.88647461 C102.49536781 51.88314369 102.49536781 51.88314369 103.90562439 51.87974548 C106 52 106 52 107 53 C107.09340434 54.62674778 107.11745171 56.25754051 107.11352539 57.88696289 C107.11340454 58.94258423 107.11328369 59.99820557 107.11315918 61.08581543 C107.10804321 62.2034729 107.10292725 63.32113037 107.09765625 64.47265625 C107.09664917 65.49387573 107.09564209 66.51509521 107.09460449 67.56726074 C107.08935415 71.39901851 107.07539303 75.23076033 107.0625 79.0625 C107.041875 87.621875 107.02125 96.18125 107 105 C89.84 105.33 72.68 105.66 55 106 C54.67 123.16 54.34 140.32 54 158 C36.18 158 18.36 158 0 158 C-0.020625 149.440625 -0.04125 140.88125 -0.0625 132.0625 C-0.071604 129.35683838 -0.08070801 126.65117676 -0.09008789 123.86352539 C-0.09300685 121.73323618 -0.09555545 119.60294642 -0.09765625 117.47265625 C-0.10277222 116.35499878 -0.10788818 115.23734131 -0.11315918 114.08581543 C-0.11334045 112.50238342 -0.11334045 112.50238342 -0.11352539 110.88696289 C-0.115746 109.96540909 -0.11796661 109.04385529 -0.12025452 108.09437561 C0 106 0 106 1 105 C2.65738443 104.90653085 4.31874644 104.88255023 5.97875977 104.88647461 C7.03978409 104.88655014 8.10080841 104.88662567 9.19398499 104.88670349 C10.348134 104.89186478 11.50228302 104.89702606 12.69140625 104.90234375 C13.86638168 104.9037587 15.04135712 104.90517365 16.25193787 104.90663147 C20.02215064 104.91225008 23.79230504 104.92480574 27.5625 104.9375 C30.11132727 104.9425126 32.66015547 104.94707592 35.20898438 104.95117188 C41.47269709 104.96137669 47.73628284 104.98094848 54 105 C54 87.84 54 70.68 54 53 C36.18 53 18.36 53 0 53 C0 70.16 0 87.32 0 105 C-18.15 105 -36.3 105 -55 105 C-55 87.51 -55 70.02 -55 52 C-28.27 51.505 -28.27 51.505 -1 51 C-0.67 34.17 -0.34 17.34 0 0 Z " fill="#FEFEFE" transform="translate(55,653)"/>
<path d="M0 0 C53.13 0 106.26 0 161 0 C161 17.49 161 34.98 161 53 C143.51 53 126.02 53 108 53 C108 70.49 108 87.98 108 106 C90.18 106 72.36 106 54 106 C54 88.51 54 71.02 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F7F7F7" transform="translate(594,0)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 52.14 54 104.28 54 158 C36.18 158 18.36 158 0 158 C0 140.51 0 123.02 0 105 C-17.39735426 105.03961002 -17.39735426 105.03961002 -34.79467773 105.09008789 C-36.96598258 105.09300684 -39.13728796 105.09555545 -41.30859375 105.09765625 C-42.44784302 105.10277222 -43.58709229 105.10788818 -44.76086426 105.11315918 C-45.83678833 105.11328003 -46.9127124 105.11340088 -48.02124023 105.11352539 C-48.96055893 105.115746 -49.89987762 105.11796661 -50.86766052 105.12025452 C-53 105 -53 105 -54 104 C-54.09340434 102.37325222 -54.11745171 100.74245949 -54.11352539 99.11303711 C-54.11340454 98.05741577 -54.11328369 97.00179443 -54.11315918 95.91418457 C-54.10548523 94.23769836 -54.10548523 94.23769836 -54.09765625 92.52734375 C-54.09664917 91.50612427 -54.09564209 90.48490479 -54.09460449 89.43273926 C-54.08935415 85.60098149 -54.07539303 81.76923967 -54.0625 77.9375 C-54.0315625 65.0984375 -54.0315625 65.0984375 -54 52 C-36.18 52 -18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(970,495)"/>
<path d="M0 0 C0 3.58679852 -0.72413825 4.34595861 -2.8125 7.1875 C-5.10140555 10.34683442 -7.36057229 13.51379 -9.52734375 16.7578125 C-15.50564165 25.68446113 -21.89226468 33.94826859 -29 42 C-29.66 42.75925781 -30.32 43.51851562 -31 44.30078125 C-32.12638558 45.59562182 -33.25753577 46.88634092 -34.39453125 48.171875 C-35.50950067 49.44147521 -36.61013736 50.72374914 -37.69921875 52.015625 C-41.16716857 56.09923332 -44.77297164 59.71264173 -48.86328125 63.171875 C-51.13655621 65.1168342 -53.31075649 67.14860655 -55.5 69.1875 C-66.40991678 78.99641601 -78.44554246 87.33533388 -91.03515625 94.82958984 C-92.31799823 95.59374795 -93.59686542 96.36462995 -94.87109375 97.14306641 C-128.51661518 117.65580899 -168.43914086 128.48669904 -207.72705078 128.20581055 C-210.39234893 128.18738003 -213.05730047 128.18530293 -215.72265625 128.18554688 C-217.44791963 128.18063539 -219.17318069 128.17480868 -220.8984375 128.16796875 C-221.67988129 128.16685593 -222.46132507 128.1657431 -223.26644897 128.16459656 C-236.90225666 128.04887167 -236.90225666 128.04887167 -241 126 C-240.55352497 121.15272752 -238.5666557 119.05628215 -235.19238281 115.65893555 C-234.69308258 115.15101974 -234.19378235 114.64310394 -233.67935181 114.11979675 C-232.03066168 112.44845518 -230.36770399 110.79222562 -228.703125 109.13671875 C-227.55016527 107.97852379 -226.39772705 106.81980946 -225.24578857 105.66059875 C-222.83127853 103.23568651 -220.40943534 100.81840151 -217.98242188 98.40600586 C-214.87216628 95.31295368 -211.78274084 92.19999621 -208.69871902 89.08081341 C-206.32435499 86.68449873 -203.9384206 84.29997661 -201.54891205 81.91877174 C-200.40482179 80.77550197 -199.26457457 79.628373 -198.12827301 78.47736168 C-196.538961 76.87064394 -194.93454829 75.28070096 -193.32519531 73.6940918 C-192.41554016 72.78539841 -191.50588501 71.87670502 -190.56866455 70.94047546 C-188 69 -188 69 -185.27931213 68.63452148 C-183 69 -183 69 -181.20581055 70.15356445 C-179.5383473 72.7069203 -179.65885733 74.5080118 -179.70703125 77.54296875 C-179.7215332 79.15268555 -179.7215332 79.15268555 -179.73632812 80.79492188 C-179.76146484 81.91447266 -179.78660156 83.03402344 -179.8125 84.1875 C-179.83280273 85.88422852 -179.83280273 85.88422852 -179.85351562 87.61523438 C-179.88890042 90.41063317 -179.93827052 93.20507892 -180 96 C-143.53250316 88.25829676 -109.75293558 68.97157126 -88.65234375 37.59375 C-83.40003038 29.34898386 -78.84149486 20.99299257 -75 12 C-72.14447237 13.2979671 -70.11891706 14.69873873 -67.875 16.875 C-59.47036503 24.31546689 -48.78707553 25.65488546 -38 25 C-26.04562108 23.10881379 -17.02236391 15.35876895 -8.4609375 7.3125 C-5.73011391 4.74639275 -2.90929666 2.35888918 0 0 Z " fill="#B32969" transform="translate(716,511)"/>
<path d="M0 0 C-0.33 17.49 -0.66 34.98 -1 53 C-18.82 53 -36.64 53 -55 53 C-55.020625 44.79125 -55.04125 36.5825 -55.0625 28.125 C-55.071604 25.53285645 -55.08070801 22.94071289 -55.09008789 20.27001953 C-55.09300744 18.22428438 -55.0955559 16.17854865 -55.09765625 14.1328125 C-55.10277222 13.06345459 -55.10788818 11.99409668 -55.11315918 10.89233398 C-55.11328003 9.87743896 -55.11340088 8.86254395 -55.11352539 7.81689453 C-55.115746 6.93309113 -55.11796661 6.04928772 -55.12025452 5.13870239 C-55 3 -55 3 -54 1 C-35.98006074 -0.14802798 -18.05409976 -0.07429671 0 0 Z M-110 53 C-91.85 53 -73.7 53 -55 53 C-54.3374034 56.97557962 -53.87591624 60.08900959 -53.88647461 63.99560547 C-53.88659546 64.94910889 -53.88671631 65.9026123 -53.88684082 66.88500977 C-53.89195679 67.86912842 -53.89707275 68.85324707 -53.90234375 69.8671875 C-53.90335083 70.78508057 -53.90435791 71.70297363 -53.90539551 72.64868164 C-53.91060341 76.05746725 -53.9245646 79.46623496 -53.9375 82.875 C-53.9684375 94.321875 -53.9684375 94.321875 -54 106 C-36.51 106 -19.02 106 -1 106 C-1 123.49 -1 140.98 -1 159 C-14.0865625 159.0309375 -14.0865625 159.0309375 -27.4375 159.0625 C-30.19536865 159.071604 -32.9532373 159.08070801 -35.79467773 159.09008789 C-37.96598258 159.09300684 -40.13728796 159.09555545 -42.30859375 159.09765625 C-43.44784302 159.10277222 -44.58709229 159.10788818 -45.76086426 159.11315918 C-46.83678833 159.11328003 -47.9127124 159.11340088 -49.02124023 159.11352539 C-49.96055893 159.115746 -50.89987762 159.11796661 -51.86766052 159.12025452 C-54 159 -54 159 -55 158 C-55.09340434 156.37325222 -55.11745171 154.74245949 -55.11352539 153.11303711 C-55.11340454 152.05741577 -55.11328369 151.00179443 -55.11315918 149.91418457 C-55.10804321 148.7965271 -55.10292725 147.67886963 -55.09765625 146.52734375 C-55.09664917 145.50612427 -55.09564209 144.48490479 -55.09460449 143.43273926 C-55.08935415 139.60098149 -55.07539303 135.76923967 -55.0625 131.9375 C-55.041875 123.378125 -55.02125 114.81875 -55 106 C-72.82 106 -90.64 106 -109 106 C-109.33 88.51 -109.66 71.02 -110 53 Z " fill="#FEFEFE" transform="translate(864,705)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.51 53.33 19.02 53.66 1 54 C0.67 71.16 0.34 88.32 0 106 C-17.49 106.33 -34.98 106.66 -53 107 C-53.33 123.83 -53.66 140.66 -54 158 C-71.49 158 -88.98 158 -107 158 C-107 140.84 -107 123.68 -107 106 C-89.51 105.67 -72.02 105.34 -54 105 C-54.03960937 88.26084826 -54.03960937 88.26084826 -54.09008789 71.52172852 C-54.09300686 69.43245494 -54.09555546 67.34318081 -54.09765625 65.25390625 C-54.10277222 64.15784058 -54.10788818 63.0617749 -54.11315918 61.93249512 C-54.11334045 60.37951721 -54.11334045 60.37951721 -54.11352539 58.79516602 C-54.115746 57.89137711 -54.11796661 56.9875882 -54.12025452 56.05641174 C-54 54 -54 54 -53 53 C-51.34261557 52.90653085 -49.68125356 52.88255023 -48.02124023 52.88647461 C-46.94531616 52.88659546 -45.86939209 52.88671631 -44.76086426 52.88684082 C-43.05199036 52.89451477 -43.05199036 52.89451477 -41.30859375 52.90234375 C-39.74727722 52.90385437 -39.74727722 52.90385437 -38.15441895 52.90539551 C-34.24876816 52.91064599 -30.34313303 52.92460711 -26.4375 52.9375 C-17.713125 52.958125 -8.98875 52.97875 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(970,53)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.92234436 0.00684998 4.99826843 0.00697083 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C33.15453552 0.07837952 41.87891052 0.09900452 50.86766052 0.12025452 C50.86766052 34.77025452 50.86766052 69.42025452 50.86766052 105.12025452 C15.22766052 105.12025452 -20.41233948 105.12025452 -57.13233948 105.12025452 C-57.13233948 54.12025452 -57.13233948 54.12025452 -56.13233948 53.12025452 C-54.47495504 53.02678536 -52.81359304 53.00280474 -51.15357971 53.00672913 C-50.09255539 53.00680466 -49.03153107 53.00688019 -47.93835449 53.00695801 C-46.78420547 53.01211929 -45.63005646 53.01728058 -44.44093323 53.02259827 C-43.26595779 53.02401321 -42.09098236 53.02542816 -40.88040161 53.02688599 C-37.11018884 53.0325046 -33.34003444 53.04506026 -29.56983948 53.05775452 C-27.02101221 53.06276712 -24.47218401 53.06733044 -21.9233551 53.07142639 C-15.65966315 53.08248007 -9.39600548 53.0992363 -3.13233948 53.12025452 C-3.13456009 52.47101517 -3.1367807 51.82177582 -3.1390686 51.15286255 C-3.16111949 44.42137703 -3.17624525 37.6899017 -3.18727112 30.95838928 C-3.19231311 28.44308557 -3.1991465 25.9277848 -3.20777893 23.41249084 C-3.21985042 19.80595677 -3.22556897 16.19946129 -3.22999573 12.59291077 C-3.23515701 11.46063553 -3.2403183 10.32836029 -3.24563599 9.16177368 C-3.24571152 8.12077011 -3.24578705 7.07976654 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#FEFEFE" transform="translate(973.1323394775391,105.87974548339844)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.90744461 0.00680466 4.96846893 0.00688019 6.06164551 0.00695801 C7.79286903 0.01469994 7.79286903 0.01469994 9.55906677 0.02259827 C10.73404221 0.02401321 11.90901764 0.02542816 13.11959839 0.02688599 C16.88981116 0.0325046 20.65996556 0.04506026 24.43016052 0.05775452 C26.97898779 0.06276712 29.52781599 0.06733044 32.0766449 0.07142639 C38.34035761 0.0816312 44.60394336 0.10120299 50.86766052 0.12025452 C51.19766052 17.28025452 51.52766052 34.44025452 51.86766052 52.12025452 C69.35766052 52.45025452 86.84766052 52.78025452 104.86766052 53.12025452 C104.86766052 70.28025452 104.86766052 87.44025452 104.86766052 105.12025452 C87.04766052 105.12025452 69.22766052 105.12025452 50.86766052 105.12025452 C50.86766052 87.96025452 50.86766052 70.80025452 50.86766052 53.12025452 C33.37766052 53.45025452 15.88766052 53.78025452 -2.13233948 54.12025452 C-2.46233948 70.95025452 -2.79233948 87.78025452 -3.13233948 105.12025452 C-20.62233948 105.12025452 -38.11233948 105.12025452 -56.13233948 105.12025452 C-56.13233948 87.96025452 -56.13233948 70.80025452 -56.13233948 53.12025452 C-38.64233948 53.12025452 -21.15233948 53.12025452 -3.13233948 53.12025452 C-3.17194918 36.05200152 -3.17194918 36.05200152 -3.22242737 18.98377991 C-3.22534633 16.8534907 -3.22789493 14.72320094 -3.22999573 12.59291077 C-3.23511169 11.4752533 -3.24022766 10.35759583 -3.24549866 9.20606995 C-3.24567993 7.62263794 -3.24567993 7.62263794 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#FEFEFE" transform="translate(435.13233947753906,105.87974548339844)"/>
<path d="M0 0 C1.43904694 0.00102722 1.43904694 0.00102722 2.90716553 0.0020752 C5.67782087 0.00859285 8.44817633 0.02500396 11.21875 0.046875 C12.05024567 0.05126587 12.88174133 0.05565674 13.73843384 0.06018066 C18.41999014 0.11649906 22.88077823 0.47909978 27.5 1.25 C28.17669678 3.02304077 28.17669678 3.02304077 28.5 5.25 C27.409729 7.04263306 27.409729 7.04263306 25.67285156 8.88134766 C25.02094849 9.57947571 24.36904541 10.27760376 23.6973877 10.99688721 C22.97224976 11.74041443 22.24711182 12.48394165 21.5 13.25 C20.76100464 14.01431335 20.02200928 14.77862671 19.26062012 15.56610107 C16.77002205 18.11221302 14.25579922 20.63285866 11.734375 23.1484375 C10.81916077 24.06460846 9.90394653 24.98077942 8.96099854 25.92471313 C7.03974333 27.8474303 5.11672231 29.76835817 3.19238281 31.68798828 C0.72880501 34.14582921 -1.73020086 36.60818799 -4.18793106 39.07187462 C-6.5447369 41.43315876 -8.9053404 43.7906306 -11.265625 46.1484375 C-12.14688049 47.03171722 -13.02813599 47.91499695 -13.93609619 48.82504272 C-14.75414734 49.63994171 -15.57219849 50.4548407 -16.41503906 51.29443359 C-17.13338928 52.01198822 -17.8517395 52.72954285 -18.59185791 53.46884155 C-21.49079696 56.17486109 -23.05102733 57.21061643 -27.0625 57.5625 C-28.196875 57.459375 -29.33125 57.35625 -30.5 57.25 C-32.73413013 53.89880481 -32.73847762 52.8322245 -32.6953125 48.92578125 C-32.68564453 47.38374023 -32.68564453 47.38374023 -32.67578125 45.81054688 C-32.65064453 44.20276367 -32.65064453 44.20276367 -32.625 42.5625 C-32.61597656 41.47904297 -32.60695313 40.39558594 -32.59765625 39.27929688 C-32.5740734 36.6026429 -32.54116126 33.92643203 -32.5 31.25 C-68.10229911 38.255082 -99.50644976 55.96227547 -120.5 86.25 C-127.10895162 96.14119005 -132.90061183 106.26580716 -137.5 117.25 C-138.44875 116.38375 -139.3975 115.5175 -140.375 114.625 C-150.0010328 106.40195174 -159.15395632 102.64964714 -171.87109375 102.87890625 C-183.04662145 104.02172125 -192.04950479 110.486606 -199.609375 118.48046875 C-201.5 120.25 -201.5 120.25 -204.25 120.5 C-204.9925 120.4175 -205.735 120.335 -206.5 120.25 C-204.89777213 115.15471635 -201.80130845 111.40047995 -198.5625 107.25 C-197.69286621 106.12440674 -197.69286621 106.12440674 -196.80566406 104.97607422 C-192.36758053 99.27014014 -187.77122214 93.71878561 -183.0546875 88.2421875 C-180.60314638 85.37081059 -178.23440595 82.44721643 -175.875 79.5 C-169.47513732 71.65132705 -162.25681976 64.74065108 -154.5 58.25 C-153.68233154 57.56164062 -153.68233154 57.56164062 -152.84814453 56.859375 C-121.58790838 30.63951052 -85.97424859 10.77609098 -45.5 3.25 C-44.75282715 3.10191895 -44.0056543 2.95383789 -43.23583984 2.80126953 C-28.89599978 0.06861078 -14.54410998 -0.01511265 0 0 Z " fill="#12A17D" transform="translate(518.5,313.75)"/>
<path d="M0 0 C4 0 4 0 5.9375 1.8125 C6.618125 2.534375 7.29875 3.25625 8 4 C8.9075 4.53625 9.815 5.0725 10.75 5.625 C11.4925 6.07875 12.235 6.5325 13 7 C13 7.66 13 8.32 13 9 C14.0828125 9.0928125 14.0828125 9.0928125 15.1875 9.1875 C18.88222728 10.25486566 20.32884822 12.25793269 23 15 C24.70859799 16.46188799 26.43842601 17.89928955 28.1875 19.3125 C29.14269531 20.08722656 30.09789062 20.86195313 31.08203125 21.66015625 C32.9702346 23.17425773 34.86317329 24.68248072 36.76171875 26.18359375 C43.29642512 31.35079804 48.87158772 36.81097466 54.3203125 43.1015625 C55.62149629 44.57220278 56.98650043 45.98650043 58.375 47.375 C73.41221672 62.41221672 86.33399184 80.04853519 96 99 C96.30115723 99.5779834 96.60231445 100.1559668 96.91259766 100.75146484 C104.30994548 114.95393125 110.8339891 129.49974081 115 145 C115.19835449 145.7204248 115.39670898 146.44084961 115.60107422 147.18310547 C123.23536616 175.29879834 123.42214238 203.09948336 123 232 C117.61441947 231.6263271 114.92781039 229.65412552 111.27001953 225.93286133 C110.73269699 225.40590668 110.19537445 224.87895203 109.64176941 224.33602905 C107.87590144 222.59718235 106.12897283 220.84065168 104.3828125 219.08203125 C103.15893138 217.86406008 101.9343831 216.64675895 100.709198 215.43009949 C98.14737626 212.88014933 95.59505138 210.32113799 93.04882812 207.75561523 C89.78542879 204.46931235 86.49781626 201.20851845 83.20245552 197.9543047 C80.66961595 195.44703939 78.15100617 192.9258546 75.63637924 190.40033531 C74.42965998 189.19212942 73.21834094 187.98849952 72.00238419 186.78959084 C70.30462633 185.11179815 68.62718671 183.41598263 66.95361328 181.71411133 C66.44874893 181.22296341 65.94388458 180.73181549 65.42372131 180.2257843 C62.99963392 177.71909575 62.03549212 176.26395532 61.56539917 172.76786804 C62 170 62 170 64 168 C66.43017578 167.77294922 66.43017578 167.77294922 69.4453125 167.8046875 C71.05986328 167.81435547 71.05986328 167.81435547 72.70703125 167.82421875 C73.83496094 167.84097656 74.96289062 167.85773438 76.125 167.875 C77.26066406 167.88402344 78.39632812 167.89304687 79.56640625 167.90234375 C82.37781299 167.92596902 85.18880298 167.95890987 88 168 C83.58956696 148.17733086 75.71760425 129.93023947 63 114 C62.57235352 113.4548877 62.14470703 112.90977539 61.70410156 112.34814453 C54.42269641 103.1371927 46.55933299 95.79229225 37 89 C36.08879395 88.34257812 36.08879395 88.34257812 35.15917969 87.671875 C26.23968819 81.28403486 17.07771345 76.31697796 7 72 C8.18883856 68.67575948 9.33065668 66.37648852 11.8125 63.875 C19.36061531 55.17704894 20.93571908 46.43455472 20.41015625 35.2421875 C19.38844226 22.25873562 10.72463821 12.12029034 1.46875 3.55859375 C0 2 0 2 0 0 Z " fill="#B5296A" transform="translate(553,279)"/>
<path d="M0 0 C2.61181641 -0.35375977 2.61181641 -0.35375977 6 0 C8.34080607 1.82730611 10.19972124 3.52061729 12.2109375 5.66015625 C12.78276764 6.24284775 13.35459778 6.82553925 13.9437561 7.42588806 C15.76885647 9.29109864 17.57228223 11.17567147 19.375 13.0625 C21.75274361 15.51666652 24.13834747 17.96313229 26.5234375 20.41015625 C27.09275497 20.99774719 27.66207245 21.58533813 28.24864197 22.19073486 C31.81800036 25.85730146 35.47099553 29.34026577 39.41772461 32.60473633 C41.6896484 34.60813772 43.58133336 36.87415915 45.48046875 39.2265625 C48.32148228 42.54229551 51.46200285 45.51781812 54.7109375 48.4296875 C55.59007812 49.23664063 56.46921875 50.04359375 57.375 50.875 C58.26960938 51.67679687 59.16421875 52.47859375 60.0859375 53.3046875 C62 56 62 56 61.9140625 59.7578125 C61.61242187 60.82773437 61.31078125 61.89765625 61 63 C58.44276771 64.27861615 56.63262898 64.11336609 53.7734375 64.09765625 C52.2265625 64.09282227 52.2265625 64.09282227 50.6484375 64.08789062 C49.56820312 64.07951172 48.48796875 64.07113281 47.375 64.0625 C45.74304688 64.05573242 45.74304688 64.05573242 44.078125 64.04882812 C41.38536211 64.03701776 38.69270812 64.02054778 36 64 C42.32332591 95.73445549 59.61317907 123.36923361 86.38671875 142.07421875 C95.72932816 148.23636538 105.98605359 153.03997646 116 158 C116 162.69475512 115.46939999 162.96226471 112.3125 166.125 C103.91480387 175.14805648 101.5374923 184.18801335 101.6640625 196.30078125 C102.72486832 207.98198023 109.82700401 217.05544179 118 225 C117.67 225.99 117.34 226.98 117 228 C112.7497269 225.97606043 108.79313929 223.79969805 105 221 C105 220.34 105 219.68 105 219 C104.38125 218.690625 103.7625 218.38125 103.125 218.0625 C101.75 217.375 100.375 216.6875 99 216 C99 215.34 99 214.68 99 214 C98.34 214 97.68 214 97 214 C97 213.34 97 212.68 97 212 C96.46375 211.938125 95.9275 211.87625 95.375 211.8125 C91.82973843 210.59964736 89.7407608 208.55389074 87 206 C87 205.34 87 204.68 87 204 C86.41863281 203.73445312 85.83726562 203.46890625 85.23828125 203.1953125 C79.01533013 199.87206112 74.23816846 194.31692071 69.7421875 188.9921875 C67.40406647 186.31855135 64.86519856 183.88359424 62.28515625 181.4453125 C61 180 61 180 61 178 C60.34 178 59.68 178 59 178 C57.28412987 176.05965224 55.69760817 174.11529177 54.125 172.0625 C53.6403125 171.43496826 53.155625 170.80743652 52.65625 170.16088867 C31.14959882 142.08161188 13.09422512 111.02726636 6 76 C5.82871582 75.154375 5.65743164 74.30875 5.48095703 73.4375 C0.72404059 49.1922933 -0.4740763 24.66290776 0 0 Z " fill="#6F2A6E" transform="translate(346,443)"/>
<path d="M0 0 C3.06722177 0.28133354 3.93666526 0.92587954 5.97265625 3.30859375 C6.66230469 4.34113281 7.35195313 5.37367188 8.0625 6.4375 C8.44680176 7.01242187 8.83110352 7.58734375 9.22705078 8.1796875 C10.50293746 10.10855494 11.75425044 12.05154407 13 14 C13.4326416 14.67305176 13.8652832 15.34610352 14.31103516 16.03955078 C49.22881354 70.74961072 49.22881354 70.74961072 43.27734375 98.3515625 C39.86902882 109.25265073 34.03058199 118.72298377 24.09765625 124.765625 C11.85745724 131.12497177 0.13138221 133.20251392 -13.33984375 129.03515625 C-25.33061871 124.3691425 -33.45267178 116.56798348 -38.8125 104.9453125 C-44.86237185 89.94003824 -41.72307127 74.65991396 -35.72412109 60.14208984 C-26.42132208 38.72799872 -14.47983735 18.31918816 0 0 Z " fill="#EFBFC9" transform="translate(510,410)"/>
<path d="M0 0 C8.435625 -0.268125 16.87125 -0.53625 25.5625 -0.8125 C28.1929126 -0.93085205 30.8233252 -1.0492041 33.53344727 -1.17114258 C44.51699675 -1.45793805 53.44241301 -1.62599197 61.8515625 6.15625 C64.03104041 8.34123988 66.02113056 10.63410653 68 13 C69.03619717 14.13243963 70.07813784 15.25965516 71.1262207 16.38110352 C83.95438876 30.37981421 93.18478894 47.60356212 98.9375 65.625 C99.14930908 66.28822266 99.36111816 66.95144531 99.5793457 67.63476562 C100.65636013 71.2141063 101.08625146 74.28204551 101 78 C100.27820557 78.02505615 99.55641113 78.0501123 98.81274414 78.07592773 C95.562465 78.19151302 92.31250312 78.31440774 89.0625 78.4375 C87.92619141 78.47681641 86.78988281 78.51613281 85.61914062 78.55664062 C84.53955078 78.59853516 83.45996094 78.64042969 82.34765625 78.68359375 C81.34742432 78.72025146 80.34719238 78.75690918 79.31665039 78.79467773 C77.03930812 78.74671841 77.03930812 78.74671841 76 80 C75.32742158 82.72091557 75.32742158 82.72091557 76 86 C78.00661531 88.83556287 80.48372804 91.13323272 83 93.515625 C83.71027344 94.21266541 84.42054688 94.90970581 85.15234375 95.62786865 C87.42114906 97.84988484 89.70929947 100.05058158 92 102.25 C94.28709717 104.46706441 96.56989732 106.68832106 98.84765625 108.91497803 C100.26592299 110.29917966 101.69028474 111.67716774 103.12109375 113.04840088 C103.76175781 113.66954773 104.40242187 114.29069458 105.0625 114.93066406 C105.63097656 115.47660217 106.19945312 116.02254028 106.78515625 116.58502197 C108 118 108 118 108 120 C107.34 120 106.68 120 106 120 C105.67 121.98 105.34 123.96 105 126 C88.17 126 71.34 126 54 126 C54 101.91 54 77.82 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FAFAFA" transform="translate(540,369)"/>
<path d="M0 0 C1.01452744 -0.00637985 2.02905487 -0.0127597 3.07432556 -0.01933289 C4.17845291 -0.02044571 5.28258026 -0.02155853 6.42016602 -0.02270508 C8.10892601 -0.02769768 8.10892601 -0.02769768 9.83180237 -0.03279114 C12.21843048 -0.03786527 14.60506572 -0.04019931 16.99169922 -0.04003906 C20.65482201 -0.04222484 24.31764349 -0.06037373 27.98071289 -0.0793457 C30.2938629 -0.08227958 32.60701434 -0.08426442 34.92016602 -0.08520508 C36.02226913 -0.09239059 37.12437225 -0.09957611 38.25987244 -0.10697937 C39.78639183 -0.10236443 39.78639183 -0.10236443 41.34375 -0.09765625 C42.24230209 -0.09908127 43.14085419 -0.10050629 44.06663513 -0.10197449 C46.23657227 0.14526367 46.23657227 0.14526367 48.23657227 2.14526367 C48.46362305 4.20825195 48.46362305 4.20825195 48.43188477 6.71557617 C48.42543945 7.61147461 48.41899414 8.50737305 48.41235352 9.43041992 C48.3955957 10.36756836 48.37883789 11.3047168 48.36157227 12.27026367 C48.35254883 13.21514648 48.34352539 14.1600293 48.33422852 15.13354492 C48.31061749 17.47103659 48.27768743 19.80802491 48.23657227 22.14526367 C49.2292234 22.14193275 49.2292234 22.14193275 50.2419281 22.13853455 C57.10317446 22.11648402 63.96441083 22.10135805 70.82568359 22.09033203 C73.38948983 22.08528997 75.95329318 22.07845653 78.51708984 22.06982422 C82.19312248 22.05775303 85.86911724 22.05203425 89.54516602 22.04760742 C90.69931503 22.04244614 91.85346405 22.03728485 93.04258728 22.03196716 C94.63412376 22.03185387 94.63412376 22.03185387 96.2578125 22.03173828 C97.1971312 22.02951767 98.13644989 22.02729706 99.10423279 22.02500916 C101.23657227 22.14526367 101.23657227 22.14526367 102.23657227 23.14526367 C102.33504193 24.70525415 102.36455844 26.26966912 102.3659668 27.83276367 C102.36911896 28.83049805 102.37227112 29.82823242 102.3755188 30.85620117 C102.37248245 32.48428711 102.37248245 32.48428711 102.36938477 34.14526367 C102.37034149 35.2512793 102.37129822 36.35729492 102.37228394 37.49682617 C102.37296593 39.84057675 102.37111031 42.1843292 102.36694336 44.52807617 C102.3615954 48.12968155 102.36688773 51.73116221 102.37329102 55.33276367 C102.37263024 57.60359728 102.37134908 59.87443081 102.36938477 62.14526367 C102.371409 63.2306543 102.37343323 64.31604492 102.3755188 65.43432617 C102.37079056 66.93092773 102.37079056 66.93092773 102.3659668 68.45776367 C102.3651712 69.34077148 102.36437561 70.2237793 102.36355591 71.13354492 C102.23657227 73.14526367 102.23657227 73.14526367 101.23657227 74.14526367 C99.61078009 74.26808319 97.97980223 74.32308871 96.34960938 74.35058594 C95.3086058 74.37053116 94.26760223 74.39047638 93.1950531 74.411026 C92.06277786 74.42773849 90.93050262 74.44445099 89.76391602 74.46166992 C88.61113663 74.48245102 87.45835724 74.50323212 86.27064514 74.52464294 C82.5718507 74.59026331 78.87298267 74.64908122 75.17407227 74.70776367 C72.67341348 74.75093702 70.17276225 74.79455091 67.67211914 74.83862305 C61.52701565 74.94595735 55.38183823 75.0477001 49.23657227 75.14526367 C48.09511219 80.69414075 48.01672537 86.15265179 47.92016602 91.79370117 C47.90151489 92.69193604 47.88286377 93.5901709 47.86364746 94.515625 C47.79567964 97.85041064 47.73532115 101.18534787 47.67407227 104.52026367 C47.52969727 111.98651367 47.38532227 119.45276367 47.23657227 127.14526367 C29.74657227 127.14526367 12.25657227 127.14526367 -5.76342773 127.14526367 C-5.78405273 118.58588867 -5.80467773 110.02651367 -5.82592773 101.20776367 C-5.83503174 98.50210205 -5.84413574 95.79644043 -5.85351562 93.00878906 C-5.85643459 90.87849985 -5.85898319 88.74821009 -5.86108398 86.61791992 C-5.86619995 85.50026245 -5.87131592 84.38260498 -5.87658691 83.2310791 C-5.87670776 82.17545776 -5.87682861 81.11983643 -5.87695312 80.03222656 C-5.87917374 79.11067276 -5.88139435 78.18911896 -5.88368225 77.23963928 C-5.76342773 75.14526367 -5.76342773 75.14526367 -4.76342773 74.14526367 C-3.13667996 74.05185933 -1.50588722 74.02781196 0.12353516 74.03173828 C1.70696716 74.03191956 1.70696716 74.03191956 3.3223877 74.03210449 C4.9988739 74.03977844 4.9988739 74.03977844 6.70922852 74.04760742 C8.24105774 74.04911804 8.24105774 74.04911804 9.80383301 74.05065918 C13.63559077 74.05590952 17.46733259 74.06987064 21.29907227 74.08276367 C29.85844727 74.10338867 38.41782227 74.12401367 47.23657227 74.14526367 C47.23657227 56.98526367 47.23657227 39.82526367 47.23657227 22.14526367 C40.63657227 22.14526367 34.03657227 22.14526367 27.23657227 22.14526367 C21.31787774 22.0041023 15.4030427 21.84621058 9.48657227 21.64526367 C7.98788382 21.59679296 6.48918585 21.54861549 4.99047852 21.50073242 C1.40572814 21.38558816 -2.17888089 21.26659871 -5.76342773 21.14526367 C-5.7923092 17.8327818 -5.81018573 14.520332 -5.82592773 11.20776367 C-5.83430664 10.26223633 -5.84268555 9.31670898 -5.85131836 8.3425293 C-5.85454102 7.4434082 -5.85776367 6.54428711 -5.86108398 5.61791992 C-5.8663208 4.78526611 -5.87155762 3.9526123 -5.87695312 3.09472656 C-5.65231376 -0.76279033 -3.3125194 0.01406468 0 0 Z " fill="#EFEFEF" transform="translate(114.763427734375,472.854736328125)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55 17.49 55 34.98 55 53 C37.18 53.33 19.36 53.66 1 54 C0.67 71.16 0.34 88.32 0 106 C-17.49 106 -34.98 106 -53 106 C-53 88.51 -53 71.02 -53 53 C-35.51 53 -18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(324,53)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.51 52.33 19.02 52.66 1 53 C0.67 70.16 0.34 87.32 0 105 C-18.15 105 -36.3 105 -55 105 C-55 87.51 -55 70.02 -55 52 C-36.85 52 -18.7 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(55,706)"/>
<path d="M0 0 C0.9215538 0.00222061 1.8431076 0.00444122 2.79258728 0.00672913 C3.83359085 0.00680466 4.87459442 0.00688019 5.94714355 0.00695801 C7.07941879 0.01211929 8.21169403 0.01728058 9.37828064 0.02259827 C11.10744972 0.02472069 11.10744972 0.02472069 12.87155151 0.02688599 C16.57043503 0.03250446 20.26925903 0.0450601 23.96812439 0.05775452 C26.46877456 0.06276714 28.96942567 0.06733045 31.47007751 0.07142639 C37.61528027 0.0824799 43.76044808 0.099236 49.90562439 0.12025452 C51.0941123 2.49723033 51.03244135 3.94668261 51.03501892 6.59828186 C51.03817108 7.52619537 51.04132324 8.45410889 51.04457092 9.41014099 C51.04153458 10.91793625 51.04153458 10.91793625 51.03843689 12.45619202 C51.03939362 13.48708954 51.04035034 14.51798706 51.04133606 15.5801239 C51.04201749 17.76407431 51.04016577 19.94802673 51.03599548 22.13197327 C51.03065759 25.47446762 51.03593613 28.81682693 51.04234314 32.15931702 C51.04168214 34.27910898 51.04040052 36.39890086 51.03843689 38.51869202 C51.04046112 39.51984039 51.04248535 40.52098877 51.04457092 41.55247498 C51.03984268 42.95380173 51.03984268 42.95380173 51.03501892 44.38343811 C51.03422333 45.20347321 51.03342773 46.0235083 51.03260803 46.86839294 C50.90562439 49.12025452 50.90562439 49.12025452 49.90562439 53.12025452 C32.41562439 53.45025452 14.92562439 53.78025452 -3.09437561 54.12025452 C-3.05484425 69.36282608 -3.05484425 69.36282608 -3.00428772 84.60536194 C-3.00136628 86.52048181 -2.99881826 88.43560231 -2.99671936 90.35072327 C-2.99160339 91.33995789 -2.98648743 92.3291925 -2.98121643 93.34840393 C-2.98103516 94.77884033 -2.98103516 94.77884033 -2.98085022 96.23817444 C-2.97862961 97.06202133 -2.976409 97.88586823 -2.97412109 98.73468018 C-3.09437561 101.12025452 -3.09437561 101.12025452 -4.09437561 106.12025452 C-21.58437561 106.12025452 -39.07437561 106.12025452 -57.09437561 106.12025452 C-57.09437561 88.63025452 -57.09437561 71.14025452 -57.09437561 53.12025452 C-39.60437561 53.12025452 -22.11437561 53.12025452 -4.09437561 53.12025452 C-4.09437561 45.86025452 -4.09437561 38.60025452 -4.09437561 31.12025452 C-3.97921489 25.67829771 -3.84597249 20.24640642 -3.65687561 14.80775452 C-3.61696546 13.47117183 -3.57725225 12.13458325 -3.53773499 10.79798889 C-3.47489319 8.92143616 -3.47489319 8.92143616 -3.41078186 7.00697327 C-3.37412415 5.89539856 -3.33746643 4.78382385 -3.29969788 3.63856506 C-3.01716378 0.17323902 -3.01716378 0.17323902 0 0 Z " fill="#F2F2F2" transform="translate(328.09437561035156,863.8797454833984)"/>
<path d="M0 0 C1.58669495 -0.00472824 1.58669495 -0.00472824 3.20544434 -0.009552 C4.93196228 -0.00651566 4.93196228 -0.00651566 6.69335938 -0.00341797 C8.45226501 -0.00485306 8.45226501 -0.00485306 10.2467041 -0.00631714 C12.73169 -0.00699917 15.21667766 -0.00514331 17.70166016 -0.00097656 C21.52054825 0.00437134 25.33931872 -0.00092083 29.15820312 -0.00732422 C31.56575547 -0.00666344 33.97330774 -0.00538229 36.38085938 -0.00341797 C37.53187134 -0.0054422 38.6828833 -0.00746643 39.86877441 -0.009552 C40.92657104 -0.00639984 41.98436768 -0.00324768 43.07421875 0 C44.47867249 0.00119339 44.47867249 0.00119339 45.91149902 0.00241089 C48.03710938 0.12939453 48.03710938 0.12939453 49.03710938 1.12939453 C49.13044643 2.72550435 49.1545631 4.32572881 49.15063477 5.92456055 C49.15051392 6.95987915 49.15039307 7.99519775 49.15026855 9.06188965 C49.14515259 10.15795532 49.14003662 11.254021 49.13476562 12.38330078 C49.13375854 13.38486206 49.13275146 14.38642334 49.13171387 15.41833496 C49.12646367 19.17619972 49.11250255 22.93404822 49.09960938 26.69189453 C49.07898438 35.08626953 49.05835938 43.48064453 49.03710938 52.12939453 C31.21710938 52.12939453 13.39710938 52.12939453 -4.96289062 52.12939453 C-4.96289062 57.40939453 -4.96289062 62.68939453 -4.96289062 68.12939453 C-5.00953085 71.26538723 -5.06278777 74.39708574 -5.14648438 77.53173828 C-5.17622093 78.69280846 -5.17622093 78.69280846 -5.20655823 79.87733459 C-5.24829945 81.47237117 -5.29116851 83.06737866 -5.33520508 84.66235352 C-5.40174238 87.11675744 -5.46066739 89.57128027 -5.51953125 92.02587891 C-5.56138996 93.59034438 -5.6036899 95.15479813 -5.64648438 96.71923828 C-5.66319687 97.45134018 -5.67990936 98.18344208 -5.6971283 98.93772888 C-5.8484929 104.01499681 -5.8484929 104.01499681 -6.96289062 105.12939453 C-8.55352372 105.22793876 -10.1485054 105.25738147 -11.7421875 105.25878906 C-13.26882019 105.2635173 -13.26882019 105.2635173 -14.82629395 105.26834106 C-15.93355835 105.26631683 -17.04082275 105.2642926 -18.18164062 105.26220703 C-19.30985229 105.26316376 -20.43806396 105.26412048 -21.60046387 105.2651062 C-23.99129288 105.26578821 -26.38212374 105.2639325 -28.77294922 105.25976562 C-32.44698214 105.25441769 -36.12089279 105.25970996 -39.79492188 105.26611328 C-42.1113284 105.2654525 -44.42773484 105.26417135 -46.74414062 105.26220703 C-47.85140503 105.26423126 -48.95866943 105.26625549 -50.0994873 105.26834106 C-51.11724243 105.2651889 -52.13499756 105.26203674 -53.18359375 105.25878906 C-54.08436646 105.25799347 -54.98513916 105.25719788 -55.91320801 105.25637817 C-57.96289062 105.12939453 -57.96289062 105.12939453 -58.96289062 104.12939453 C-59.06143485 102.53876143 -59.09087756 100.94377976 -59.09228516 99.35009766 C-59.09543732 98.33234253 -59.09858948 97.3145874 -59.10183716 96.26599121 C-59.09981293 95.15872681 -59.0977887 94.0514624 -59.09570312 92.91064453 C-59.09665985 91.78243286 -59.09761658 90.65422119 -59.09860229 89.49182129 C-59.0992843 87.10099227 -59.0974286 84.71016142 -59.09326172 82.31933594 C-59.08791378 78.64530302 -59.09320605 74.97139236 -59.09960938 71.29736328 C-59.0989486 68.98095676 -59.09766744 66.66455031 -59.09570312 64.34814453 C-59.09873947 62.68724792 -59.09873947 62.68724792 -59.10183716 60.99279785 C-59.098685 59.97504272 -59.09553284 58.9572876 -59.09228516 57.90869141 C-59.09148956 57.0079187 -59.09069397 56.107146 -59.08987427 55.17907715 C-58.96289062 53.12939453 -58.96289062 53.12939453 -57.96289062 52.12939453 C-56.33614285 52.03599019 -54.70535011 52.01194282 -53.07592773 52.01586914 C-52.03492416 52.01594467 -50.99392059 52.0160202 -49.92137146 52.01609802 C-48.78909622 52.02125931 -47.65682098 52.02642059 -46.49023438 52.03173828 C-45.33745499 52.03315323 -44.1846756 52.03456818 -42.9969635 52.036026 C-39.29807999 52.04164448 -35.59925598 52.05420012 -31.90039062 52.06689453 C-29.39974045 52.07190715 -26.89908934 52.07647047 -24.3984375 52.08056641 C-18.25323474 52.09161991 -12.10806693 52.10837601 -5.96289062 52.12939453 C-5.96511124 51.49268326 -5.96733185 50.85597198 -5.96961975 50.19996643 C-5.99167103 43.59824177 -6.00679656 36.99652749 -6.01782227 30.39477539 C-6.02286419 27.9279742 -6.02969753 25.46117601 -6.03833008 22.99438477 C-6.05040187 19.45734924 -6.05612018 15.92035308 -6.06054688 12.38330078 C-6.06570816 11.27289932 -6.07086945 10.16249786 -6.07618713 9.01844788 C-6.07626266 7.99746506 -6.0763382 6.97648224 -6.07641602 5.92456055 C-6.07863663 5.02077164 -6.08085724 4.11698273 -6.08314514 3.18580627 C-5.84796921 -0.83581861 -3.47102337 0.00294939 0 0 Z " fill="#F0F0F0" transform="translate(167.962890625,316.87060546875)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.51 53.33 19.02 53.66 1 54 C0.67 71.16 0.34 88.32 0 106 C-17.49 106 -34.98 106 -53 106 C-53 88.51 -53 71.02 -53 53 C-35.51 53 -18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(916,211)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.92234436 0.00684998 4.99826843 0.00697083 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C33.15453552 0.07837952 41.87891052 0.09900452 50.86766052 0.12025452 C50.86766052 17.61025452 50.86766052 35.10025452 50.86766052 53.12025452 C33.37766052 53.45025452 15.88766052 53.78025452 -2.13233948 54.12025452 C-2.09273011 70.85940626 -2.09273011 70.85940626 -2.04225159 87.598526 C-2.03933262 89.68779957 -2.03678401 91.77707371 -2.03468323 93.86634827 C-2.02956726 94.96241394 -2.02445129 96.05847961 -2.0191803 97.1877594 C-2.01899902 98.7407373 -2.01899902 98.7407373 -2.01881409 100.3250885 C-2.01659348 101.22887741 -2.01437286 102.13266632 -2.01208496 103.06384277 C-2.13233948 105.12025452 -2.13233948 105.12025452 -3.13233948 106.12025452 C-4.78972391 106.21372367 -6.45108592 106.23770429 -8.11109924 106.23377991 C-9.18702332 106.23365906 -10.26294739 106.23353821 -11.37147522 106.2334137 C-12.51072449 106.22829773 -13.64997375 106.22318176 -14.82374573 106.21791077 C-16.38506226 106.21640015 -16.38506226 106.21640015 -17.97792053 106.21485901 C-21.88357131 106.20960852 -25.78920645 106.19564741 -29.69483948 106.18275452 C-38.41921448 106.16212952 -47.14358948 106.14150452 -56.13233948 106.12025452 C-56.13233948 88.63025452 -56.13233948 71.14025452 -56.13233948 53.12025452 C-38.64233948 53.12025452 -21.15233948 53.12025452 -3.13233948 53.12025452 C-3.17194918 36.05200152 -3.17194918 36.05200152 -3.22242737 18.98377991 C-3.22534633 16.8534907 -3.22789493 14.72320094 -3.22999573 12.59291077 C-3.23511169 11.4752533 -3.24022766 10.35759583 -3.24549866 9.20606995 C-3.24567993 7.62263794 -3.24567993 7.62263794 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#FEFEFE" transform="translate(919.1323394775391,52.87974548339844)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.51 53.33 19.02 53.66 1 54 C0.67 71.16 0.34 88.32 0 106 C-17.49 106 -34.98 106 -53 106 C-53 88.51 -53 71.02 -53 53 C-35.51 53 -18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0F0" transform="translate(432,53)"/>
<path d="M0 0 C1.1821995 0.00138269 1.1821995 0.00138269 2.38828182 0.00279331 C3.28997097 0.00141865 4.19166012 0.00004398 5.12067318 -0.00137234 C6.6160738 0.00402058 6.6160738 0.00402058 8.14168453 0.00952244 C9.18546261 0.00937641 10.22924068 0.00923038 11.3046484 0.00907993 C14.77305295 0.00977956 18.24140454 0.0175743 21.70979977 0.02539158 C24.1073367 0.02725558 26.50487401 0.02867957 28.90241146 0.0296793 C35.22684936 0.03350589 41.55126446 0.04333737 47.87569332 0.05438328 C55.45640498 0.06638823 63.03712424 0.07099897 70.61784267 0.07683659 C82.14720883 0.08654905 93.67652492 0.10570464 105.20589352 0.12304783 C104.87589352 17.61304783 104.54589352 35.10304783 104.20589352 53.12304783 C68.89589352 53.12304783 33.58589352 53.12304783 -2.79410648 53.12304783 C-2.79410648 0.19163229 -2.79410648 0.19163229 0 0 Z " fill="#F2F2F2" transform="translate(381.7941064834595,810.8769521713257)"/>
<path d="M0 0 C0.95708359 0.00222061 1.91416718 0.00444122 2.9002533 0.00672913 C3.98129837 0.00680466 5.06234344 0.00688019 6.17614746 0.00695801 C7.94018166 0.01469994 7.94018166 0.01469994 9.73985291 0.02259827 C10.93702438 0.02401321 12.13419586 0.02542816 13.36764526 0.02688599 C17.20918732 0.03250472 21.05067208 0.04506041 24.89219666 0.05775452 C27.48920102 0.0627671 30.0862063 0.06733043 32.68321228 0.07142639 C39.06541382 0.08163138 45.44749076 0.10120316 51.82969666 0.12025452 C51.82969666 17.61025452 51.82969666 35.10025452 51.82969666 53.12025452 C34.00969666 53.45025452 16.18969666 53.78025452 -2.17030334 54.12025452 C-2.50030334 70.95025452 -2.83030334 87.78025452 -3.17030334 105.12025452 C-20.66030334 105.12025452 -38.15030334 105.12025452 -56.17030334 105.12025452 C-56.17030334 87.96025452 -56.17030334 70.80025452 -56.17030334 53.12025452 C-38.68030334 53.12025452 -21.19030334 53.12025452 -3.17030334 53.12025452 C-3.20991305 36.05200152 -3.20991305 36.05200152 -3.26039124 18.98377991 C-3.2633102 16.8534907 -3.2658588 14.72320094 -3.26795959 12.59291077 C-3.27307556 11.4752533 -3.27819153 10.35759583 -3.28346252 9.20606995 C-3.2836438 7.62263794 -3.2836438 7.62263794 -3.28382874 6.00721741 C-3.28604935 5.0856636 -3.28826996 4.1641098 -3.29055786 3.21463013 C-3.12491431 0.32975042 -2.88616406 0.1599197 0 0 Z " fill="#FEFEFE" transform="translate(327.17030334472656,105.87974548339844)"/>
<path d="M0 0 C0.95708359 0.00222061 1.91416718 0.00444122 2.9002533 0.00672913 C3.98129837 0.00680466 5.06234344 0.00688019 6.17614746 0.00695801 C7.94018166 0.01469994 7.94018166 0.01469994 9.73985291 0.02259827 C10.93702438 0.02401321 12.13419586 0.02542816 13.36764526 0.02688599 C17.20918732 0.03250472 21.05067208 0.04506041 24.89219666 0.05775452 C27.48920102 0.0627671 30.0862063 0.06733043 32.68321228 0.07142639 C39.06541382 0.08163138 45.44749076 0.10120316 51.82969666 0.12025452 C51.82969666 17.28025452 51.82969666 34.44025452 51.82969666 52.12025452 C34.00969666 52.45025452 16.18969666 52.78025452 -2.17030334 53.12025452 C-2.50030334 70.28025452 -2.83030334 87.44025452 -3.17030334 105.12025452 C-20.66030334 105.12025452 -38.15030334 105.12025452 -56.17030334 105.12025452 C-56.17030334 87.63025452 -56.17030334 70.14025452 -56.17030334 52.12025452 C-38.68030334 52.12025452 -21.19030334 52.12025452 -3.17030334 52.12025452 C-3.20991271 35.38110278 -3.20991271 35.38110278 -3.26039124 18.64198303 C-3.26331021 16.55270946 -3.26585881 14.46343532 -3.26795959 12.37416077 C-3.27307556 11.27809509 -3.27819153 10.18202942 -3.28346252 9.05274963 C-3.2836438 7.49977173 -3.2836438 7.49977173 -3.28382874 5.91542053 C-3.28604935 5.01163162 -3.28826996 4.10784271 -3.29055786 3.17666626 C-3.12334243 0.3171997 -2.86095594 0.15852294 0 0 Z " fill="#EFEFEF" transform="translate(327.17030334472656,158.87974548339844)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55 17.49 55 34.98 55 53 C72.82 53 90.64 53 109 53 C109 69.83 109 86.66 109 104 C91.18 104 73.36 104 55 104 C54.67 87.5 54.34 71 54 54 C50.26945312 53.93941406 46.53890625 53.87882812 42.6953125 53.81640625 C39.09454242 53.75465285 35.49380491 53.69125023 31.89306641 53.62768555 C29.38463216 53.58429097 26.87616751 53.5426193 24.36767578 53.50268555 C20.76846132 53.44509243 17.16940058 53.38136657 13.5703125 53.31640625 C12.44319855 53.29969376 11.31608459 53.28298126 10.15481567 53.26576233 C9.11388763 53.24581711 8.07295959 53.22587189 7.00048828 53.20532227 C6.08115509 53.18977798 5.1618219 53.1742337 4.21463013 53.15821838 C2 53 2 53 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFF0EF" transform="translate(0,369)"/>
<path d="M0 0 C1.37899979 0.00666183 1.37899979 0.00666183 2.78585815 0.01345825 C4.36910889 0.0138208 4.36910889 0.0138208 5.98434448 0.01419067 C7.09688599 0.02442261 8.20942749 0.03465454 9.35568237 0.04519653 C10.37589478 0.04721069 11.39610718 0.04922485 12.44723511 0.05130005 C16.26832558 0.06178587 20.08935212 0.08970832 23.91036987 0.11550903 C32.44911987 0.15675903 40.98786987 0.19800903 49.78536987 0.24050903 C49.78536987 17.73050903 49.78536987 35.22050903 49.78536987 53.24050903 C31.96536987 53.24050903 14.14536987 53.24050903 -4.21463013 53.24050903 C-4.25588013 44.86675903 -4.29713013 36.49300903 -4.33963013 27.86550903 C-4.35783813 25.22115845 -4.37604614 22.57680786 -4.39480591 19.85232544 C-4.40064496 17.76557621 -4.4057419 15.67882471 -4.40994263 13.59207153 C-4.42017456 12.50112183 -4.43040649 11.41017212 -4.44094849 10.28616333 C-4.44119019 9.25096558 -4.44143188 8.21576782 -4.44168091 7.14920044 C-4.44612213 6.24763214 -4.45056335 5.34606384 -4.45513916 4.41717529 C-4.11038039 1.29702312 -3.11276564 0.33804663 0 0 Z M-54.12025452 53.12025452 C-53.19870071 53.12247513 -52.27714691 53.12469574 -51.32766724 53.12698364 C-49.74423523 53.12716492 -49.74423523 53.12716492 -48.1288147 53.12734985 C-46.45232849 53.1350238 -46.45232849 53.1350238 -44.74197388 53.14285278 C-43.21014465 53.1443634 -43.21014465 53.1443634 -41.64736938 53.14590454 C-37.81561162 53.15115488 -33.9838698 53.165116 -30.15213013 53.17800903 C-21.59275513 53.19863403 -13.03338013 53.21925903 -4.21463013 53.24050903 C-4.21463013 70.73050903 -4.21463013 88.22050903 -4.21463013 106.24050903 C-21.70463013 106.24050903 -39.19463013 106.24050903 -57.21463013 106.24050903 C-57.23525513 97.68113403 -57.25588013 89.12175903 -57.27713013 80.30300903 C-57.28623413 77.59734741 -57.29533813 74.89168579 -57.30471802 72.10403442 C-57.30763698 69.97374522 -57.31018558 67.84345545 -57.31228638 65.71316528 C-57.31740234 64.59550781 -57.32251831 63.47785034 -57.32778931 62.32632446 C-57.32791016 61.27070312 -57.32803101 60.21508179 -57.32815552 59.12747192 C-57.33037613 58.20591812 -57.33259674 57.28436432 -57.33488464 56.33488464 C-57.17203251 53.49862073 -56.95651843 53.28310665 -54.12025452 53.12025452 Z " fill="#FEFEFE" transform="translate(920.2146301269531,810.7594909667969)"/>
<path d="M0 0 C0.92042587 0.02009628 1.84085175 0.04019257 2.78916931 0.06089783 C3.75923416 0.08793289 4.72929901 0.11496796 5.72875977 0.14282227 C6.7398732 0.16643326 7.75098663 0.19004425 8.79273987 0.21437073 C12.00204107 0.29055477 15.21107291 0.37477237 18.42016602 0.45922852 C20.60439791 0.51249457 22.78864269 0.56523461 24.97290039 0.61743164 C30.30965328 0.74610815 35.64620828 0.88136982 40.98266602 1.02172852 C42.16044682 6.5886786 42.11027349 12.01087415 42.08032227 17.67016602 C42.07890732 18.6826944 42.07749237 19.69522278 42.07603455 20.73843384 C42.07045745 23.95789602 42.05790914 27.17728751 42.04516602 30.39672852 C42.04014806 32.58552959 42.03558567 34.77433176 42.03149414 36.96313477 C42.02049552 42.31602329 42.00378022 47.66887085 41.98266602 53.02172852 C35.09588067 53.16486402 28.20907907 53.3071972 21.32226562 53.44897461 C18.97981389 53.49729264 16.63736593 53.54579383 14.29492188 53.59448242 C10.92652344 53.66446399 7.55811197 53.73378527 4.18969727 53.80297852 C2.62068413 53.83578918 2.62068413 53.83578918 1.01997375 53.8692627 C0.03933456 53.88928345 -0.94130463 53.9093042 -1.95166016 53.92993164 C-3.24072517 53.95657898 -3.24072517 53.95657898 -4.55583191 53.98376465 C-7.0427357 54.02212029 -9.53013443 54.02172852 -12.01733398 54.02172852 C-12.01733398 71.18172852 -12.01733398 88.34172852 -12.01733398 106.02172852 C-29.83733398 106.02172852 -47.65733398 106.02172852 -66.01733398 106.02172852 C-66.03795898 97.46235352 -66.05858398 88.90297852 -66.07983398 80.08422852 C-66.08893799 77.37856689 -66.09804199 74.67290527 -66.10742188 71.88525391 C-66.11034084 69.7549647 -66.11288944 67.62467494 -66.11499023 65.49438477 C-66.1201062 64.37672729 -66.12522217 63.25906982 -66.13049316 62.10754395 C-66.13061401 61.05192261 -66.13073486 59.99630127 -66.13085938 58.90869141 C-66.13307999 57.9871376 -66.1353006 57.0655838 -66.1375885 56.11610413 C-66.01733398 54.02172852 -66.01733398 54.02172852 -65.01733398 53.02172852 C-63.35994955 52.92825936 -61.69858755 52.90427874 -60.03857422 52.90820312 C-58.9775499 52.90827866 -57.91652557 52.90835419 -56.823349 52.90843201 C-55.66919998 52.91359329 -54.51505096 52.91875458 -53.32592773 52.92407227 C-52.1509523 52.92548721 -50.97597687 52.92690216 -49.76539612 52.92835999 C-45.99518335 52.9339786 -42.22502895 52.94653426 -38.45483398 52.95922852 C-35.90600671 52.96424112 -33.35717852 52.96880444 -30.80834961 52.97290039 C-24.54463689 52.9831052 -18.28105114 53.00267699 -12.01733398 53.02172852 C-12.01733398 35.86172852 -12.01733398 18.70172852 -12.01733398 1.02172852 C-4.14233398 -0.10327148 -4.14233398 -0.10327148 0 0 Z " fill="#EDEDED" transform="translate(660.017333984375,704.978271484375)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.90744461 0.00680466 4.96846893 0.00688019 6.06164551 0.00695801 C7.79286903 0.01469994 7.79286903 0.01469994 9.55906677 0.02259827 C10.73404221 0.02401321 11.90901764 0.02542816 13.11959839 0.02688599 C16.88981116 0.0325046 20.65996556 0.04506026 24.43016052 0.05775452 C26.97898779 0.06276712 29.52781599 0.06733044 32.0766449 0.07142639 C38.34035761 0.0816312 44.60394336 0.10120299 50.86766052 0.12025452 C50.86766052 17.28025452 50.86766052 34.44025452 50.86766052 52.12025452 C33.37766052 52.12025452 15.88766052 52.12025452 -2.13233948 52.12025452 C-2.42172547 69.18840444 -2.42172547 69.18840444 -2.70045471 86.25672913 C-2.73855912 88.38702582 -2.77702665 90.51731607 -2.81593323 92.64759827 C-2.83240906 93.76525574 -2.84888489 94.88291321 -2.86585999 96.03443909 C-2.88604187 97.09006042 -2.90622375 98.14568176 -2.92701721 99.23329163 C-2.94256149 100.15484543 -2.95810577 101.07639923 -2.97412109 102.02587891 C-3.13233948 104.12025452 -3.13233948 104.12025452 -4.13233948 105.12025452 C-5.72297258 105.21879874 -7.31795425 105.24824145 -8.91163635 105.24964905 C-10.43826904 105.25437729 -10.43826904 105.25437729 -11.9957428 105.25920105 C-13.1030072 105.25717682 -14.21027161 105.25515259 -15.35108948 105.25306702 C-16.47930115 105.25402374 -17.60751282 105.25498047 -18.76991272 105.25596619 C-21.16074174 105.25664819 -23.55157259 105.25479249 -25.94239807 105.25062561 C-29.61643099 105.24527767 -33.29034164 105.25056994 -36.96437073 105.25697327 C-39.28077725 105.25631249 -41.59718369 105.25503133 -43.91358948 105.25306702 C-45.02085388 105.25509125 -46.12811829 105.25711548 -47.26893616 105.25920105 C-48.28669128 105.25604889 -49.30444641 105.25289673 -50.3530426 105.24964905 C-51.25381531 105.24885345 -52.15458801 105.24805786 -53.08265686 105.24723816 C-55.13233948 105.12025452 -55.13233948 105.12025452 -56.13233948 104.12025452 C-56.22574382 102.49350674 -56.24979119 100.862714 -56.24586487 99.23329163 C-56.24574402 98.17767029 -56.24562317 97.12204895 -56.24549866 96.03443909 C-56.23782471 94.35795288 -56.23782471 94.35795288 -56.22999573 92.64759827 C-56.22898865 91.62637878 -56.22798157 90.6051593 -56.22694397 89.55299377 C-56.22169363 85.72123601 -56.20773251 81.88949419 -56.19483948 78.05775452 C-56.16390198 65.21869202 -56.16390198 65.21869202 -56.13233948 52.12025452 C-38.64233948 52.12025452 -21.15233948 52.12025452 -3.13233948 52.12025452 C-3.17194885 35.38110278 -3.17194885 35.38110278 -3.22242737 18.64198303 C-3.22534634 16.55270946 -3.22789494 14.46343532 -3.22999573 12.37416077 C-3.23511169 11.27809509 -3.24022766 10.18202942 -3.24549866 9.05274963 C-3.24567993 7.49977173 -3.24567993 7.49977173 -3.24586487 5.91542053 C-3.24808548 5.01163162 -3.25030609 4.10784271 -3.25259399 3.17666626 C-3.08677921 0.34115132 -2.8362359 0.15995116 0 0 Z " fill="#F0F0F0" transform="translate(919.1323394775391,316.87974548339844)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C4.4603064 0.0069104 4.4603064 0.0069104 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C37.51672302 0.08869202 37.51672302 0.08869202 50.86766052 0.12025452 C50.86766052 24.21025452 50.86766052 48.30025452 50.86766052 73.12025452 C42.32891052 73.16150452 33.79016052 73.20275452 24.99266052 73.24525452 C20.9478241 73.27256653 20.9478241 73.27256653 16.8212738 73.3004303 C14.69350891 73.3062693 12.56574179 73.31136626 10.43797302 73.31556702 C9.32543152 73.32579895 8.21289001 73.33603088 7.06663513 73.34657288 C5.4833844 73.34693542 5.4833844 73.34693542 3.8681488 73.3473053 C2.94881561 73.35174652 2.02948242 73.35618774 1.08229065 73.36076355 C-1.13233948 73.12025452 -1.13233948 73.12025452 -3.13233948 71.12025452 C-3.37957764 68.22900391 -3.37957764 68.22900391 -3.3752594 64.48329163 C-3.37715775 63.80185593 -3.37905609 63.12042023 -3.38101196 62.41833496 C-3.38472293 60.16130646 -3.37401217 57.90459826 -3.36280823 55.64759827 C-3.36161661 54.08343544 -3.36116323 52.5192719 -3.36141968 50.95510864 C-3.35985432 47.67572048 -3.35155999 44.39644141 -3.33815002 41.11708069 C-3.32114607 36.9044778 -3.31733604 32.69199472 -3.31809521 28.47936153 C-3.31782387 25.24956103 -3.31234877 22.01978694 -3.30509377 18.78999519 C-3.30190229 17.23618838 -3.29993858 15.68237856 -3.29920006 14.12856865 C-3.29704232 11.96160101 -3.28831095 9.79476289 -3.27760315 7.62782288 C-3.27379135 6.39253342 -3.26997955 5.15724396 -3.26605225 3.88452148 C-3.08657071 0.17406894 -3.08657071 0.17406894 0 0 Z " fill="#EFF0EF" transform="translate(919.1323394775391,421.87974548339844)"/>
<path d="M0 0 C15.51 0 31.02 0 47 0 C47.04010881 17.92863777 47.04010881 17.92863777 47.04882812 25.54492188 C47.0548162 30.75090549 47.06191555 35.95687159 47.07543945 41.1628418 C47.08626959 45.35790258 47.0922771 49.55294459 47.09487724 53.74801826 C47.09673126 55.35206968 47.10035144 56.95612003 47.10573006 58.5601635 C47.11294219 60.79916515 47.11399087 63.0380883 47.11352539 65.27709961 C47.115746 66.55395126 47.11796661 67.83080292 47.12025452 69.14634705 C47 72 47 72 46 73 C42.89748799 73.08874135 39.8173188 73.11518455 36.71484375 73.09765625 C35.78402481 73.0962413 34.85320587 73.09482635 33.8941803 73.09336853 C30.90858809 73.08775172 27.92306971 73.0751964 24.9375 73.0625 C22.91862087 73.05748716 20.89974057 73.05292388 18.88085938 73.04882812 C13.92054428 73.03777683 8.96028468 73.02050095 4 73 C3.98018066 72.07477539 3.96036133 71.14955078 3.93994141 70.19628906 C4.51941379 42.71570248 4.51941379 42.71570248 0 16 C0 10.72 0 5.44 0 0 Z " fill="#FEFEFE" transform="translate(763,422)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55 17.82 55 35.64 55 54 C36.85 54 18.7 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#EFEFEF" transform="translate(0,970)"/>
<path d="M0 0 C3.98580921 3.54366398 7.12882011 7.58330744 10.25 11.875 C10.96506714 12.85738647 10.96506714 12.85738647 11.69458008 13.85961914 C19.65424311 24.95382214 26.14662277 36.73768969 32.05029297 49.03125 C32.97853189 50.95549644 33.92706099 52.8685939 34.87890625 54.78125 C43.63038805 72.62044983 49.72689894 92.25566618 44.03125 112.05859375 C39.43285363 125.17447432 32.08982873 134.30059334 20.1484375 141.4921875 C6.1582889 148.19218422 -9.32889796 148.87879251 -24 144 C-36.77840132 138.57395847 -46.60113152 130.16958748 -52.15234375 117.3359375 C-54.27659516 111.84765807 -55.62137283 106.86872111 -56 101 C-56.0515625 100.36320312 -56.103125 99.72640625 -56.15625 99.0703125 C-57.19469881 76.13790122 -44.91377801 51.83356141 -33 33 C-32.01865827 31.33461309 -31.03953381 29.66791788 -30.0625 28 C-26.94784816 22.81967233 -23.54471731 17.89371903 -20 13 C-19.23945313 11.93523437 -18.47890625 10.87046875 -17.6953125 9.7734375 C-16.90203489 8.68156936 -16.10777697 7.59041273 -15.3125 6.5 C-14.58675781 5.4996875 -13.86101562 4.499375 -13.11328125 3.46875 C-9.05903686 -1.26744678 -6.00540801 -1.58037053 0 0 Z M-6 8 C-7.75080536 9.93659226 -9.24057749 11.82039506 -10.75 13.9375 C-11.22026611 14.58992676 -11.69053223 15.24235352 -12.17504883 15.91455078 C-23.02576374 31.31274773 -32.54397806 47.70128906 -40 65 C-40.73283203 66.60681641 -40.73283203 66.60681641 -41.48046875 68.24609375 C-48.00886358 82.96848562 -50.47644115 97.5626357 -45 113 C-39.71412531 124.37862745 -31.44080273 132.00286777 -20 137 C-8.68836855 141.02880024 3.0950801 139.51334731 14 135 C26.22333043 128.64386818 32.90281622 119.49875728 37.109375 106.59765625 C43.10594586 82.37466606 27.80436641 56.27977908 16 36 C12.50086664 30.22176699 8.79340553 24.58825756 5 19 C4.59797363 18.40268066 4.19594727 17.80536133 3.78173828 17.18994141 C0.61039921 12.42356511 0.61039921 12.42356511 -3 8 C-3.99 8 -4.98 8 -6 8 Z " fill="#FCF9F7" transform="translate(516,402)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.82 54 35.64 54 54 C36.18 54 18.36 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#F2F2F2" transform="translate(594,970)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.82 54 35.64 54 54 C36.18 54 18.36 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#F1F1F1" transform="translate(486,970)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.82 54 35.64 54 54 C36.18 54 18.36 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#F0F0F0" transform="translate(217,970)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.82 54 35.64 54 54 C36.18 54 18.36 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#FEFEFE" transform="translate(163,970)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.82 54 35.64 54 54 C36.18 54 18.36 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#F0F0F0" transform="translate(109,970)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.82 54 35.64 54 54 C36.18 54 18.36 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#FEFEFE" transform="translate(55,970)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55 17.49 55 34.98 55 53 C36.85 53 18.7 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(0,917)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55 17.49 55 34.98 55 53 C36.85 53 18.7 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0F0" transform="translate(0,264)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55 17.49 55 34.98 55 53 C36.85 53 18.7 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(0,0)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55.020625 8.559375 55.04125 17.11875 55.0625 25.9375 C55.071604 28.64316162 55.08070801 31.34882324 55.09008789 34.13647461 C55.09300685 36.26676382 55.09555545 38.39705358 55.09765625 40.52734375 C55.10277222 41.64500122 55.10788818 42.76265869 55.11315918 43.91418457 C55.11334045 45.49761658 55.11334045 45.49761658 55.11352539 47.11303711 C55.115746 48.03459091 55.11796661 48.95614471 55.12025452 49.90562439 C55 52 55 52 54 53 C52.31198015 53.09353163 50.62004793 53.11744791 48.92944336 53.11352539 C47.84839828 53.11344986 46.76735321 53.11337433 45.65354919 53.11329651 C43.889515 53.10555458 43.889515 53.10555458 42.08984375 53.09765625 C40.89267227 53.0962413 39.69550079 53.09482635 38.46205139 53.09336853 C34.62050934 53.08774979 30.77902457 53.07519411 26.9375 53.0625 C24.34049563 53.05748741 21.74349035 53.05292409 19.14648438 53.04882812 C12.76428284 53.03862313 6.3822059 53.01905136 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(0,53)"/>
<path d="M0 0 C8.70375 -0.04125 17.4075 -0.0825 26.375 -0.125 C29.12376465 -0.14320801 31.8725293 -0.16141602 34.70458984 -0.18017578 C36.8733704 -0.18601475 39.04215315 -0.19111171 41.2109375 -0.1953125 C42.91213745 -0.2106604 42.91213745 -0.2106604 44.64770508 -0.22631836 C46.26140991 -0.22668091 46.26140991 -0.22668091 47.90771484 -0.22705078 C48.84481293 -0.231492 49.78191101 -0.23593323 50.74740601 -0.24050903 C53 0 53 0 55 2 C55.24050903 4.17666626 55.24050903 4.17666626 55.22705078 6.90869141 C55.22680908 7.94388916 55.22656738 8.97908691 55.22631836 10.0456543 C55.21097046 11.68207886 55.21097046 11.68207886 55.1953125 13.3515625 C55.19329834 14.3521167 55.19128418 15.3526709 55.18920898 16.38354492 C55.17872374 20.13074307 55.15080129 23.87787601 55.125 27.625 C55.08375 35.99875 55.0425 44.3725 55 53 C36.85 53 18.7 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(0,864)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C-1.1497912 50.70041761 -1.12670434 49.40161935 -1.12939453 46.8449707 C-1.13254669 45.98680252 -1.13569885 45.12863434 -1.13894653 44.24446106 C-1.1369223 43.31429672 -1.13489807 42.38413239 -1.1328125 41.42578125 C-1.13376923 40.46858688 -1.13472595 39.51139252 -1.13571167 38.52519226 C-1.13639322 36.49506566 -1.13454071 34.46493689 -1.13037109 32.43481445 C-1.12505171 29.34256004 -1.13030176 26.25045282 -1.13671875 23.15820312 C-1.13605739 21.18489551 -1.13477503 19.211588 -1.1328125 17.23828125 C-1.13483673 16.31823807 -1.13686096 15.39819489 -1.13894653 14.45027161 C-1.13579437 13.57634262 -1.13264221 12.70241364 -1.12939453 11.80200195 C-1.12859894 11.04192337 -1.12780334 10.28184479 -1.12698364 9.49873352 C-0.96515789 6.31439088 -0.45091519 3.15640636 0 0 Z " fill="#EFEFEF" transform="translate(163,0)"/>
<path d="M0 0 C0.95708359 0.0199855 1.91416718 0.03997101 2.9002533 0.06056213 C3.98129837 0.08065842 5.06234344 0.1007547 6.17614746 0.12145996 C7.35217026 0.14849503 8.52819305 0.17553009 9.73985291 0.2033844 C10.93702438 0.22699539 12.13419586 0.25060638 13.36764526 0.27493286 C17.20927629 0.3517971 21.05071715 0.43572311 24.89219666 0.51979065 C27.48919241 0.57298856 30.08619758 0.62572908 32.68321228 0.67799377 C39.06552975 0.806579 45.44754146 0.94469858 51.82969666 1.08229065 C51.82969666 18.57229065 51.82969666 36.06229065 51.82969666 54.08229065 C34.00969666 54.08229065 16.18969666 54.08229065 -2.17030334 54.08229065 C-2.35592834 45.35791565 -2.54155334 36.63354065 -2.73280334 27.64479065 C-2.8247699 23.50798767 -2.8247699 23.50798767 -2.91859436 19.28761292 C-2.96253625 17.1163157 -3.00610096 14.94501081 -3.04920959 12.7736969 C-3.07591736 11.63444763 -3.10262512 10.49519836 -3.13014221 9.32142639 C-3.1505658 8.24550232 -3.17098938 7.16957825 -3.19203186 6.06105042 C-3.21201736 5.12173172 -3.23200287 4.18241302 -3.25259399 3.21463013 C-3.1400551 0.29848913 -2.91628908 0.11057594 0 0 Z " fill="#FEFEFE" transform="translate(918.1703033447266,703.9177093505859)"/>
<path d="M0 0 C0.20254517 2.21463013 0.20254517 2.21463013 0.13525391 5.00048828 C0.11470947 6.05598877 0.09416504 7.11148926 0.07299805 8.19897461 C0.02526245 9.86778687 0.02526245 9.86778687 -0.0234375 11.5703125 C-0.04510986 12.5905249 -0.06678223 13.6107373 -0.08911133 14.66186523 C-0.17328606 18.48317133 -0.27522428 22.30406942 -0.375 26.125 C-0.58125 34.66375 -0.7875 43.2025 -1 52 C-18.82 52 -36.64 52 -55 52 C-55.020625 43.440625 -55.04125 34.88125 -55.0625 26.0625 C-55.071604 23.35683838 -55.08070801 20.65117676 -55.09008789 17.86352539 C-55.09300685 15.73323618 -55.09555545 13.60294642 -55.09765625 11.47265625 C-55.10277222 10.35499878 -55.10788818 9.23734131 -55.11315918 8.08581543 C-55.11328003 7.03019409 -55.11340088 5.97457275 -55.11352539 4.88696289 C-55.115746 3.96540909 -55.11796661 3.04385529 -55.12025452 2.09437561 C-55 0 -55 0 -54 -1 C-52.38515011 -1.13322586 -50.76466175 -1.19888363 -49.14477539 -1.23706055 C-47.59295311 -1.27666145 -47.59295311 -1.27666145 -46.00978088 -1.31706238 C-44.88377975 -1.34004898 -43.75777863 -1.36303558 -42.59765625 -1.38671875 C-40.87560219 -1.42500542 -40.87560219 -1.42500542 -39.11875916 -1.46406555 C-36.68510314 -1.516181 -34.25138802 -1.56559472 -31.81762695 -1.61254883 C-28.08186463 -1.68711349 -24.34671141 -1.77773325 -20.61132812 -1.86914062 C-18.25262427 -1.91765426 -15.89390053 -1.96521226 -13.53515625 -2.01171875 C-12.41117935 -2.04077805 -11.28720245 -2.06983734 -10.12916565 -2.09977722 C-9.0914653 -2.11672134 -8.05376495 -2.13366547 -6.98461914 -2.15112305 C-6.06830215 -2.17031296 -5.15198517 -2.18950287 -4.207901 -2.20927429 C-2 -2 -2 -2 0 0 Z " fill="#FEFEFE" transform="translate(703,865)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.82 53 35.64 53 54 C35.51 54 18.02 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#F0F0F0" transform="translate(810,970)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.82 53 35.64 53 54 C35.51 54 18.02 54 0 54 C0 36.18 0 18.36 0 0 Z " fill="#F0F0F0" transform="translate(702,970)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F0F0F0" transform="translate(648,917)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F1F1F1" transform="translate(540,917)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(163,917)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(109,917)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(55,917)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(755,811)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(55,811)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(55,600)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(970,369)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(648,106)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(594,106)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(540,106)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(217,106)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(163,106)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(594,53)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(540,53)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F0F0F0" transform="translate(217,53)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(970,0)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(594,0)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(540,0)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(486,0)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(55,0)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C4.4603064 0.0069104 4.4603064 0.0069104 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C37.51672302 0.08869202 37.51672302 0.08869202 50.86766052 0.12025452 C50.86766052 17.61025452 50.86766052 35.10025452 50.86766052 53.12025452 C33.04766052 53.12025452 15.22766052 53.12025452 -3.13233948 53.12025452 C-3.15296448 44.56087952 -3.17358948 36.00150452 -3.19483948 27.18275452 C-3.20394348 24.4770929 -3.21304749 21.77143127 -3.22242737 18.98377991 C-3.22534633 16.8534907 -3.22789493 14.72320094 -3.22999573 12.59291077 C-3.23511169 11.4752533 -3.24022766 10.35759583 -3.24549866 9.20606995 C-3.24561951 8.15044861 -3.24574036 7.09482727 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#FEFEFE" transform="translate(973.1323394775391,863.8797454833984)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C4.4603064 0.0069104 4.4603064 0.0069104 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C37.51672302 0.08869202 37.51672302 0.08869202 50.86766052 0.12025452 C50.86766052 17.61025452 50.86766052 35.10025452 50.86766052 53.12025452 C33.04766052 53.12025452 15.22766052 53.12025452 -3.13233948 53.12025452 C-3.15296448 44.56087952 -3.17358948 36.00150452 -3.19483948 27.18275452 C-3.20394348 24.4770929 -3.21304749 21.77143127 -3.22242737 18.98377991 C-3.22534633 16.8534907 -3.22789493 14.72320094 -3.22999573 12.59291077 C-3.23511169 11.4752533 -3.24022766 10.35759583 -3.24549866 9.20606995 C-3.24561951 8.15044861 -3.24574036 7.09482727 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#FEFEFE" transform="translate(973.1323394775391,757.8797454833984)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C4.4603064 0.0069104 4.4603064 0.0069104 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C37.51672302 0.08869202 37.51672302 0.08869202 50.86766052 0.12025452 C50.86766052 17.61025452 50.86766052 35.10025452 50.86766052 53.12025452 C33.04766052 53.12025452 15.22766052 53.12025452 -3.13233948 53.12025452 C-3.15296448 44.56087952 -3.17358948 36.00150452 -3.19483948 27.18275452 C-3.20394348 24.4770929 -3.21304749 21.77143127 -3.22242737 18.98377991 C-3.22534633 16.8534907 -3.22789493 14.72320094 -3.22999573 12.59291077 C-3.23511169 11.4752533 -3.24022766 10.35759583 -3.24549866 9.20606995 C-3.24561951 8.15044861 -3.24574036 7.09482727 -3.24586487 6.00721741 C-3.24808548 5.0856636 -3.25030609 4.1641098 -3.25259399 3.21463013 C-3.08833702 0.35389928 -2.86123587 0.16136105 0 0 Z " fill="#FEFEFE" transform="translate(166.13233947753906,757.8797454833984)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54.020625 8.559375 54.04125 17.11875 54.0625 25.9375 C54.071604 28.64316162 54.08070801 31.34882324 54.09008789 34.13647461 C54.09300685 36.26676382 54.09555545 38.39705358 54.09765625 40.52734375 C54.10277222 41.64500122 54.10788818 42.76265869 54.11315918 43.91418457 C54.11334045 45.49761658 54.11334045 45.49761658 54.11352539 47.11303711 C54.115746 48.03459091 54.11796661 48.95614471 54.12025452 49.90562439 C54 52 54 52 53 53 C51.34261557 53.09346915 49.68125356 53.11744977 48.02124023 53.11352539 C46.94531616 53.11340454 45.86939209 53.11328369 44.76086426 53.11315918 C43.05199036 53.10548523 43.05199036 53.10548523 41.30859375 53.09765625 C39.74727722 53.09614563 39.74727722 53.09614563 38.15441895 53.09460449 C34.24876816 53.08935401 30.34313303 53.07539289 26.4375 53.0625 C17.713125 53.041875 8.98875 53.02125 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(163,600)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C45.275625 53.020625 36.55125 53.04125 27.5625 53.0625 C24.80463135 53.071604 22.0467627 53.08070801 19.20532227 53.09008789 C17.03401742 53.09300684 14.86271204 53.09555545 12.69140625 53.09765625 C11.55215698 53.10277222 10.41290771 53.10788818 9.23913574 53.11315918 C8.16321167 53.11328003 7.0872876 53.11340088 5.97875977 53.11352539 C5.03944107 53.115746 4.10012238 53.11796661 3.13233948 53.12025452 C1 53 1 53 0 52 C-0.09340434 50.37325222 -0.11745171 48.74245949 -0.11352539 47.11303711 C-0.11340454 46.05741577 -0.11328369 45.00179443 -0.11315918 43.91418457 C-0.10548523 42.23769836 -0.10548523 42.23769836 -0.09765625 40.52734375 C-0.09664917 39.50612427 -0.09564209 38.48490479 -0.09460449 37.43273926 C-0.08935415 33.60098149 -0.07539303 29.76923967 -0.0625 25.9375 C-0.0315625 13.0984375 -0.0315625 13.0984375 0 0 Z " fill="#EFEFEF" transform="translate(970,264)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54.020625 8.559375 54.04125 17.11875 54.0625 25.9375 C54.071604 28.64316162 54.08070801 31.34882324 54.09008789 34.13647461 C54.09300685 36.26676382 54.09555545 38.39705358 54.09765625 40.52734375 C54.10277222 41.64500122 54.10788818 42.76265869 54.11315918 43.91418457 C54.11334045 45.49761658 54.11334045 45.49761658 54.11352539 47.11303711 C54.115746 48.03459091 54.11796661 48.95614471 54.12025452 49.90562439 C54 52 54 52 53 53 C51.34261557 53.09346915 49.68125356 53.11744977 48.02124023 53.11352539 C46.94531616 53.11340454 45.86939209 53.11328369 44.76086426 53.11315918 C43.05199036 53.10548523 43.05199036 53.10548523 41.30859375 53.09765625 C39.74727722 53.09614563 39.74727722 53.09614563 38.15441895 53.09460449 C34.24876816 53.08935401 30.34313303 53.07539289 26.4375 53.0625 C17.713125 53.041875 8.98875 53.02125 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F0F0F0" transform="translate(217,264)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C45.275625 53.020625 36.55125 53.04125 27.5625 53.0625 C24.80463135 53.071604 22.0467627 53.08070801 19.20532227 53.09008789 C17.03401742 53.09300684 14.86271204 53.09555545 12.69140625 53.09765625 C11.55215698 53.10277222 10.41290771 53.10788818 9.23913574 53.11315918 C8.16321167 53.11328003 7.0872876 53.11340088 5.97875977 53.11352539 C5.03944107 53.115746 4.10012238 53.11796661 3.13233948 53.12025452 C1 53 1 53 0 52 C-0.09340434 50.37325222 -0.11745171 48.74245949 -0.11352539 47.11303711 C-0.11340454 46.05741577 -0.11328369 45.00179443 -0.11315918 43.91418457 C-0.10548523 42.23769836 -0.10548523 42.23769836 -0.09765625 40.52734375 C-0.09664917 39.50612427 -0.09564209 38.48490479 -0.09460449 37.43273926 C-0.08935415 33.60098149 -0.07539303 29.76923967 -0.0625 25.9375 C-0.0315625 13.0984375 -0.0315625 13.0984375 0 0 Z " fill="#EFEFEF" transform="translate(486,106)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C45.275625 53.020625 36.55125 53.04125 27.5625 53.0625 C24.80463135 53.071604 22.0467627 53.08070801 19.20532227 53.09008789 C17.03401742 53.09300684 14.86271204 53.09555545 12.69140625 53.09765625 C11.55215698 53.10277222 10.41290771 53.10788818 9.23913574 53.11315918 C8.16321167 53.11328003 7.0872876 53.11340088 5.97875977 53.11352539 C5.03944107 53.115746 4.10012238 53.11796661 3.13233948 53.12025452 C1 53 1 53 0 52 C-0.09340434 50.37325222 -0.11745171 48.74245949 -0.11352539 47.11303711 C-0.11340454 46.05741577 -0.11328369 45.00179443 -0.11315918 43.91418457 C-0.10548523 42.23769836 -0.10548523 42.23769836 -0.09765625 40.52734375 C-0.09664917 39.50612427 -0.09564209 38.48490479 -0.09460449 37.43273926 C-0.08935415 33.60098149 -0.07539303 29.76923967 -0.0625 25.9375 C-0.0315625 13.0984375 -0.0315625 13.0984375 0 0 Z " fill="#EFEFEF" transform="translate(55,106)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C4.4603064 0.0069104 4.4603064 0.0069104 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C37.51672302 0.08869202 37.51672302 0.08869202 50.86766052 0.12025452 C50.86766052 17.61025452 50.86766052 35.10025452 50.86766052 53.12025452 C42.14328552 53.14087952 33.41891052 53.16150452 24.43016052 53.18275452 C21.67229187 53.19185852 18.91442322 53.20096252 16.07298279 53.21034241 C13.90167795 53.21326136 11.73037256 53.21580996 9.55906677 53.21791077 C8.4198175 53.22302673 7.28056824 53.2281427 6.10679626 53.2334137 C5.03087219 53.23353455 3.95494812 53.2336554 2.84642029 53.23377991 C1.90710159 53.23600052 0.9677829 53.23822113 0 53.24050903 C-2.13233948 53.12025452 -2.13233948 53.12025452 -3.13233948 52.12025452 C-3.2308837 50.52962142 -3.26032641 48.93463974 -3.26173401 47.34095764 C-3.26488617 46.32320251 -3.26803833 45.30544739 -3.27128601 44.2568512 C-3.26926178 43.14958679 -3.26723755 42.04232239 -3.26515198 40.90150452 C-3.2661087 39.77329285 -3.26706543 38.64508118 -3.26805115 37.48268127 C-3.26873315 35.09185226 -3.26687745 32.7010214 -3.26271057 30.31019592 C-3.25736263 26.63616301 -3.26265491 22.96225235 -3.26905823 19.28822327 C-3.26839745 16.97181674 -3.26711629 14.6554103 -3.26515198 12.33900452 C-3.26818832 10.67810791 -3.26818832 10.67810791 -3.27128601 8.98365784 C-3.26813385 7.96590271 -3.26498169 6.94814758 -3.26173401 5.89955139 C-3.26093842 4.99877869 -3.26014282 4.09800598 -3.25932312 3.16993713 C-3.08400007 0.33999297 -2.831922 0.15970788 0 0 Z " fill="#EFEFEF" transform="translate(758.1323394775391,916.8797454833984)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C4.4603064 0.0069104 4.4603064 0.0069104 6.10679626 0.00709534 C7.81567017 0.01476929 7.81567017 0.01476929 9.55906677 0.02259827 C11.1203833 0.02410889 11.1203833 0.02410889 12.71324158 0.02565002 C16.61889236 0.03090051 20.52452749 0.04486163 24.43016052 0.05775452 C37.51672302 0.08869202 37.51672302 0.08869202 50.86766052 0.12025452 C50.86766052 17.61025452 50.86766052 35.10025452 50.86766052 53.12025452 C42.14328552 53.14087952 33.41891052 53.16150452 24.43016052 53.18275452 C21.67229187 53.19185852 18.91442322 53.20096252 16.07298279 53.21034241 C13.90167795 53.21326136 11.73037256 53.21580996 9.55906677 53.21791077 C8.4198175 53.22302673 7.28056824 53.2281427 6.10679626 53.2334137 C5.03087219 53.23353455 3.95494812 53.2336554 2.84642029 53.23377991 C1.90710159 53.23600052 0.9677829 53.23822113 0 53.24050903 C-2.13233948 53.12025452 -2.13233948 53.12025452 -3.13233948 52.12025452 C-3.2308837 50.52962142 -3.26032641 48.93463974 -3.26173401 47.34095764 C-3.26488617 46.32320251 -3.26803833 45.30544739 -3.27128601 44.2568512 C-3.26926178 43.14958679 -3.26723755 42.04232239 -3.26515198 40.90150452 C-3.2661087 39.77329285 -3.26706543 38.64508118 -3.26805115 37.48268127 C-3.26873315 35.09185226 -3.26687745 32.7010214 -3.26271057 30.31019592 C-3.25736263 26.63616301 -3.26265491 22.96225235 -3.26905823 19.28822327 C-3.26839745 16.97181674 -3.26711629 14.6554103 -3.26515198 12.33900452 C-3.26818832 10.67810791 -3.26818832 10.67810791 -3.27128601 8.98365784 C-3.26813385 7.96590271 -3.26498169 6.94814758 -3.26173401 5.89955139 C-3.26093842 4.99877869 -3.26014282 4.09800598 -3.25932312 3.16993713 C-3.08400007 0.33999297 -2.831922 0.15970788 0 0 Z " fill="#EFF0F0" transform="translate(758.1323394775391,263.87974548339844)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54.020625 8.559375 54.04125 17.11875 54.0625 25.9375 C54.071604 28.64316162 54.08070801 31.34882324 54.09008789 34.13647461 C54.09300685 36.26676382 54.09555545 38.39705358 54.09765625 40.52734375 C54.10277222 41.64500122 54.10788818 42.76265869 54.11315918 43.91418457 C54.11334045 45.49761658 54.11334045 45.49761658 54.11352539 47.11303711 C54.115746 48.03459091 54.11796661 48.95614471 54.12025452 49.90562439 C54 52 54 52 53 53 C51.37872577 53.09861598 49.75317632 53.12798767 48.12890625 53.12939453 C46.57224243 53.13412277 46.57224243 53.13412277 44.98413086 53.13894653 C43.29042358 53.13591019 43.29042358 53.13591019 41.5625 53.1328125 C39.83688843 53.13424759 39.83688843 53.13424759 38.07641602 53.13571167 C35.63850856 53.13639369 33.2005993 53.1345379 30.76269531 53.13037109 C27.01623482 53.12502317 23.26989423 53.13031539 19.5234375 53.13671875 C17.16145807 53.13605797 14.79947871 53.13477682 12.4375 53.1328125 C11.30836182 53.13483673 10.17922363 53.13686096 9.01586914 53.13894653 C7.45920532 53.13421829 7.45920532 53.13421829 5.87109375 53.12939453 C4.95255615 53.12859894 4.03401855 53.12780334 3.08764648 53.12698364 C1 53 1 53 0 52 C-0.09340434 50.37325222 -0.11745171 48.74245949 -0.11352539 47.11303711 C-0.11340454 46.05741577 -0.11328369 45.00179443 -0.11315918 43.91418457 C-0.10548523 42.23769836 -0.10548523 42.23769836 -0.09765625 40.52734375 C-0.09664917 39.50612427 -0.09564209 38.48490479 -0.09460449 37.43273926 C-0.08935415 33.60098149 -0.07539303 29.76923967 -0.0625 25.9375 C-0.0315625 13.0984375 -0.0315625 13.0984375 0 0 Z " fill="#EFEFEF" transform="translate(55,211)"/>
<path d="M0 0 C1.52179115 -0.00472824 1.52179115 -0.00472824 3.07432556 -0.009552 C4.73051659 -0.00651566 4.73051659 -0.00651566 6.42016602 -0.00341797 C8.10892601 -0.00485306 8.10892601 -0.00485306 9.83180237 -0.00631714 C12.21843522 -0.0069992 14.60506991 -0.00514311 16.99169922 -0.00097656 C20.65474603 0.00436634 24.31766995 -0.00091814 27.98071289 -0.00732422 C30.2938642 -0.00666334 32.60701544 -0.00538199 34.92016602 -0.00341797 C36.02226913 -0.0054422 37.12437225 -0.00746643 38.25987244 -0.009552 C39.78639183 -0.00482376 39.78639183 -0.00482376 41.34375 0 C42.24230209 0.00079559 43.14085419 0.00159119 44.06663513 0.00241089 C46.23657227 0.12939453 46.23657227 0.12939453 48.23657227 1.12939453 C48.23657227 18.28939453 48.23657227 35.44939453 48.23657227 53.12939453 C30.41657227 53.12939453 12.59657227 53.12939453 -5.76342773 53.12939453 C-5.78405273 44.57001953 -5.80467773 36.01064453 -5.82592773 27.19189453 C-5.83503174 24.48623291 -5.84413574 21.78057129 -5.85351562 18.99291992 C-5.85643459 16.86263071 -5.85898319 14.73234095 -5.86108398 12.60205078 C-5.86619995 11.48439331 -5.87131592 10.36673584 -5.87658691 9.21520996 C-5.87670776 8.15958862 -5.87682861 7.10396729 -5.87695312 6.01635742 C-5.87917374 5.09480362 -5.88139435 4.17324982 -5.88368225 3.22377014 C-5.6547518 -0.76332636 -3.46805262 0.00307339 0 0 Z " fill="#F0F0F0" transform="translate(222.763427734375,863.87060546875)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55.020625 8.394375 55.04125 16.78875 55.0625 25.4375 C55.071604 28.09095459 55.08070801 30.74440918 55.09008789 33.47827148 C55.09300686 35.56754506 55.09555546 37.65681919 55.09765625 39.74609375 C55.10277222 40.84215942 55.10788818 41.9382251 55.11315918 43.06750488 C55.11334045 44.62048279 55.11334045 44.62048279 55.11352539 46.20483398 C55.115746 47.10862289 55.11796661 48.0124118 55.12025452 48.94358826 C55 51 55 51 54 52 C52.31198015 52.09353163 50.62004793 52.11744791 48.92944336 52.11352539 C47.84839828 52.11344986 46.76735321 52.11337433 45.65354919 52.11329651 C43.889515 52.10555458 43.889515 52.10555458 42.08984375 52.09765625 C40.89267227 52.0962413 39.69550079 52.09482635 38.46205139 52.09336853 C34.62050934 52.08774979 30.77902457 52.07519411 26.9375 52.0625 C24.34049563 52.05748741 21.74349035 52.05292409 19.14648438 52.04882812 C12.76428284 52.03862313 6.3822059 52.01905136 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(0,653)"/>
<path d="M0 0 C18.15 0 36.3 0 55 0 C55.020625 8.394375 55.04125 16.78875 55.0625 25.4375 C55.071604 28.09095459 55.08070801 30.74440918 55.09008789 33.47827148 C55.09300686 35.56754506 55.09555546 37.65681919 55.09765625 39.74609375 C55.10277222 40.84215942 55.10788818 41.9382251 55.11315918 43.06750488 C55.11334045 44.62048279 55.11334045 44.62048279 55.11352539 46.20483398 C55.115746 47.10862289 55.11796661 48.0124118 55.12025452 48.94358826 C55 51 55 51 54 52 C52.31198015 52.09353163 50.62004793 52.11744791 48.92944336 52.11352539 C47.84839828 52.11344986 46.76735321 52.11337433 45.65354919 52.11329651 C43.889515 52.10555458 43.889515 52.10555458 42.08984375 52.09765625 C40.89267227 52.0962413 39.69550079 52.09482635 38.46205139 52.09336853 C34.62050934 52.08774979 30.77902457 52.07519411 26.9375 52.0625 C24.34049563 52.05748741 21.74349035 52.05292409 19.14648438 52.04882812 C12.76428284 52.03862313 6.3822059 52.01905136 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(0,159)"/>
<path d="M0 0 C1.01452744 -0.00637985 2.02905487 -0.0127597 3.07432556 -0.01933289 C4.17845291 -0.02044571 5.28258026 -0.02155853 6.42016602 -0.02270508 C8.10892601 -0.02769768 8.10892601 -0.02769768 9.83180237 -0.03279114 C12.21843048 -0.03786527 14.60506572 -0.04019931 16.99169922 -0.04003906 C20.65482201 -0.04222484 24.31764349 -0.06037373 27.98071289 -0.0793457 C30.2938629 -0.08227958 32.60701434 -0.08426442 34.92016602 -0.08520508 C36.02226913 -0.09239059 37.12437225 -0.09957611 38.25987244 -0.10697937 C39.78639183 -0.10236443 39.78639183 -0.10236443 41.34375 -0.09765625 C42.24230209 -0.09908127 43.14085419 -0.10050629 44.06663513 -0.10197449 C46.23657227 0.14526367 46.23657227 0.14526367 48.23657227 2.14526367 C48.4770813 4.32192993 48.4770813 4.32192993 48.46362305 7.05395508 C48.46338135 8.08915283 48.46313965 9.12435059 48.46289062 10.19091797 C48.44754272 11.82734253 48.44754272 11.82734253 48.43188477 13.49682617 C48.42987061 14.49738037 48.42785645 15.49793457 48.42578125 16.52880859 C48.41529601 20.27600674 48.38737356 24.02313968 48.36157227 27.77026367 C48.32032227 36.14401367 48.27907227 44.51776367 48.23657227 53.14526367 C30.41657227 53.14526367 12.59657227 53.14526367 -5.76342773 53.14526367 C-5.78405273 44.58588867 -5.80467773 36.02651367 -5.82592773 27.20776367 C-5.83503174 24.50210205 -5.84413574 21.79644043 -5.85351562 19.00878906 C-5.85643459 16.87849985 -5.85898319 14.74821009 -5.86108398 12.61791992 C-5.86619995 11.50026245 -5.87131592 10.38260498 -5.87658691 9.2310791 C-5.87670776 8.17545776 -5.87682861 7.11983643 -5.87695312 6.03222656 C-5.87917374 5.11067276 -5.88139435 4.18911896 -5.88368225 3.23963928 C-5.65494375 -0.74411408 -3.46773823 0.01472372 0 0 Z " fill="#F0F0F0" transform="translate(114.763427734375,863.854736328125)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C54.22721424 2.45442848 54.12691608 4.05717514 54.12939453 6.80102539 C54.13254669 7.79868423 54.13569885 8.79634308 54.13894653 9.82423401 C54.1369223 10.90446335 54.13489807 11.98469269 54.1328125 13.09765625 C54.13376923 14.20225693 54.13472595 15.3068576 54.13571167 16.44493103 C54.13639301 18.78270525 54.13454196 21.12048136 54.13037109 23.45825195 C54.12501716 27.05098688 54.1303203 30.64359708 54.13671875 34.23632812 C54.13605806 36.50260444 54.13477709 38.76888069 54.1328125 41.03515625 C54.13483673 42.11740982 54.13686096 43.19966339 54.13894653 44.31471252 C54.13421829 45.80647255 54.13421829 45.80647255 54.12939453 47.32836914 C54.12859894 48.20836075 54.12780334 49.08835236 54.12698364 49.99501038 C54 52 54 52 53 53 C51.34261557 53.09346915 49.68125356 53.11744977 48.02124023 53.11352539 C46.94531616 53.11340454 45.86939209 53.11328369 44.76086426 53.11315918 C43.05199036 53.10548523 43.05199036 53.10548523 41.30859375 53.09765625 C39.74727722 53.09614563 39.74727722 53.09614563 38.15441895 53.09460449 C34.24876816 53.08935401 30.34313303 53.07539289 26.4375 53.0625 C17.713125 53.041875 8.98875 53.02125 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F0F0F0" transform="translate(109,53)"/>
<path d="M0 0 C1.47095879 0.0001133 1.47095879 0.0001133 2.97163391 0.00022888 C4.54064705 0.00797081 4.54064705 0.00797081 6.14135742 0.01586914 C7.22188889 0.01728409 8.30242035 0.01869904 9.41569519 0.02015686 C12.85943393 0.02574459 16.30310715 0.0382949 19.74682617 0.05102539 C22.08471586 0.05604197 24.42260656 0.0606046 26.76049805 0.06469727 C32.4851297 0.07571001 38.20972325 0.09243598 43.93432617 0.11352539 C43.9595931 7.50080641 43.97715778 14.88807637 43.98925781 22.27539062 C43.99429981 24.79069434 44.0011332 27.30599511 44.00976562 29.82128906 C44.02183711 33.42782314 44.02755566 37.03431862 44.03198242 40.64086914 C44.03714371 41.77314438 44.04230499 42.90541962 44.04762268 44.07200623 C44.04769821 45.1130098 44.04777374 46.15401337 44.04785156 47.2265625 C44.05007217 48.1481163 44.05229279 49.0696701 44.05458069 50.01914978 C43.93432617 52.11352539 43.93432617 52.11352539 42.93432617 53.11352539 C41.27694174 53.20699454 39.61557973 53.23097516 37.95556641 53.22705078 C36.89454208 53.22697525 35.83351776 53.22689972 34.74034119 53.2268219 C33.00911766 53.21907997 33.00911766 53.21907997 31.24291992 53.21118164 C30.06794449 53.20976669 28.89296906 53.20835175 27.68238831 53.20689392 C23.91217553 53.20127531 20.14202114 53.18871965 16.37182617 53.17602539 C13.8229989 53.17101279 11.2741707 53.16644947 8.7253418 53.16235352 C2.46162908 53.15214871 -3.80195667 53.13257691 -10.06567383 53.11352539 C-10.06567383 35.95352539 -10.06567383 18.79352539 -10.06567383 1.11352539 C-6.37985054 0.37636073 -3.65443557 -0.00944299 0 0 Z " fill="#FDFDFD" transform="translate(658.065673828125,757.886474609375)"/>
<path d="M0 0 C4.455 -0.020625 8.91 -0.04125 13.5 -0.0625 C14.84771484 -0.071604 16.19542969 -0.08070801 17.58398438 -0.09008789 C29.77471266 -0.11637563 41.77225737 0.49051072 54 1 C54 18.16 54 35.32 54 53 C36.18 53 18.36 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F1F2F1" transform="translate(486,864)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.49 54 34.98 54 53 C36.51 53 19.02 53 1 53 C0.67 35.51 0.34 18.02 0 0 Z " fill="#EFEFEF" transform="translate(809,758)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 16.83 54 33.66 54 51 C49.71069382 52.71572247 48.21089419 53.24575954 43.93432617 53.13525391 C42.94009644 53.11470947 41.9458667 53.09416504 40.92150879 53.07299805 C39.37288147 53.02526245 39.37288147 53.02526245 37.79296875 52.9765625 C36.8347522 52.95489014 35.87653564 52.93321777 34.88928223 52.91088867 C31.32173236 52.82711225 27.7546329 52.72496711 24.1875 52.625 C16.205625 52.41875 8.22375 52.2125 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFF0EF" transform="translate(217,653)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(863,917)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#F0F0F0" transform="translate(271,811)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(863,758)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(863,600)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(379,53)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(271,53)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#FEFEFE" transform="translate(863,0)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(810,0)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(702,0)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(379,0)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C35.51 53 18.02 53 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFEFEF" transform="translate(271,0)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#FEFEFE" transform="translate(970,653)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#FEFEFE" transform="translate(970,548)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(55,317)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53.020625 8.559375 53.04125 17.11875 53.0625 25.9375 C53.071604 28.64316162 53.08070801 31.34882324 53.09008789 34.13647461 C53.09300685 36.26676382 53.09555545 38.39705358 53.09765625 40.52734375 C53.10277222 41.64500122 53.10788818 42.76265869 53.11315918 43.91418457 C53.11334045 45.49761658 53.11334045 45.49761658 53.11352539 47.11303711 C53.115746 48.03459091 53.11796661 48.95614471 53.12025452 49.90562439 C53 52 53 52 52 53 C50.37325222 53.09340434 48.74245949 53.11745171 47.11303711 53.11352539 C46.05741577 53.11340454 45.00179443 53.11328369 43.91418457 53.11315918 C42.23769836 53.10548523 42.23769836 53.10548523 40.52734375 53.09765625 C39.50612427 53.09664917 38.48490479 53.09564209 37.43273926 53.09460449 C33.60098149 53.08935415 29.76923967 53.07539303 25.9375 53.0625 C17.378125 53.041875 8.81875 53.02125 0 53 C0 35.51 0 18.02 0 0 Z " fill="#EFF0EF" transform="translate(109,264)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.49 53 34.98 53 53 C44.440625 53.020625 35.88125 53.04125 27.0625 53.0625 C23.00400757 53.07615601 23.00400757 53.07615601 18.86352539 53.09008789 C16.73323618 53.09300685 14.60294642 53.09555545 12.47265625 53.09765625 C11.35499878 53.10277222 10.23734131 53.10788818 9.08581543 53.11315918 C8.03019409 53.11328003 6.97457275 53.11340088 5.88696289 53.11352539 C4.50463219 53.11685631 4.50463219 53.11685631 3.09437561 53.12025452 C1 53 1 53 0 52 C-0.09340434 50.37325222 -0.11745171 48.74245949 -0.11352539 47.11303711 C-0.11340454 46.05741577 -0.11328369 45.00179443 -0.11315918 43.91418457 C-0.10548523 42.23769836 -0.10548523 42.23769836 -0.09765625 40.52734375 C-0.09664917 39.50612427 -0.09564209 38.48490479 -0.09460449 37.43273926 C-0.08935415 33.60098149 -0.07539303 29.76923967 -0.0625 25.9375 C-0.0315625 13.0984375 -0.0315625 13.0984375 0 0 Z " fill="#EFEFEF" transform="translate(810,211)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(648,159)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#FEFEFE" transform="translate(594,159)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#F0F0F0" transform="translate(540,159)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 17.16 54 34.32 54 52 C36.18 52 18.36 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(217,159)"/>
<path d="M0 0 C1.01775513 -0.00315216 2.03551025 -0.00630432 3.08410645 -0.009552 C4.19137085 -0.00752777 5.29863525 -0.00550354 6.43945312 -0.00341797 C7.56766479 -0.00437469 8.69587646 -0.00533142 9.85827637 -0.00631714 C12.24910538 -0.00699915 14.63993624 -0.00514344 17.03076172 -0.00097656 C20.70479464 0.00437137 24.37870529 -0.0009209 28.05273438 -0.00732422 C30.3691409 -0.00666344 32.68554734 -0.00538229 35.00195312 -0.00341797 C36.66284973 -0.00645432 36.66284973 -0.00645432 38.3572998 -0.009552 C39.37505493 -0.00639984 40.39281006 -0.00324768 41.44140625 0 C42.79256531 0.00119339 42.79256531 0.00119339 44.17102051 0.00241089 C46.22070312 0.12939453 46.22070312 0.12939453 47.22070312 1.12939453 C47.31410746 2.75614231 47.33815483 4.38693504 47.33422852 6.01635742 C47.33410767 7.07197876 47.33398682 8.1276001 47.3338623 9.21520996 C47.32874634 10.33286743 47.32363037 11.4505249 47.31835938 12.60205078 C47.31735229 13.62327026 47.31634521 14.64448975 47.31530762 15.69665527 C47.31005727 19.52841304 47.29609615 23.36015486 47.28320312 27.19189453 C47.26257813 35.75126953 47.24195313 44.31064453 47.22070312 53.12939453 C29.73070312 53.12939453 12.24070312 53.12939453 -5.77929688 53.12939453 C-5.79992187 44.57001953 -5.82054687 36.01064453 -5.84179688 27.19189453 C-5.85090088 24.48623291 -5.86000488 21.78057129 -5.86938477 18.99291992 C-5.87230373 16.86263071 -5.87485233 14.73234095 -5.87695312 12.60205078 C-5.88206909 11.48439331 -5.88718506 10.36673584 -5.89245605 9.21520996 C-5.8925769 8.15958862 -5.89269775 7.10396729 -5.89282227 6.01635742 C-5.89504288 5.09480362 -5.89726349 4.17324982 -5.89955139 3.22377014 C-5.67030382 -0.76884933 -3.4715873 0.00306622 0 0 Z " fill="#EFF0F0" transform="translate(707.779296875,863.87060546875)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.90744461 0.00680466 4.96846893 0.00688019 6.06164551 0.00695801 C7.21579453 0.01211929 8.36994354 0.01728058 9.55906677 0.02259827 C10.73404221 0.02401321 11.90901764 0.02542816 13.11959839 0.02688599 C16.88981116 0.0325046 20.65996556 0.04506026 24.43016052 0.05775452 C26.97898779 0.06276712 29.52781599 0.06733044 32.0766449 0.07142639 C38.34035761 0.0816312 44.60394336 0.10120299 50.86766052 0.12025452 C50.86766052 17.28025452 50.86766052 34.44025452 50.86766052 52.12025452 C33.04766052 52.12025452 15.22766052 52.12025452 -3.13233948 52.12025452 C-3.15296448 43.72587952 -3.17358948 35.33150452 -3.19483948 26.68275452 C-3.20394348 24.02929993 -3.21304749 21.37584534 -3.22242737 18.64198303 C-3.22534634 16.55270946 -3.22789494 14.46343532 -3.22999573 12.37416077 C-3.23511169 11.27809509 -3.24022766 10.18202942 -3.24549866 9.05274963 C-3.24561951 8.01743103 -3.24574036 6.98211243 -3.24586487 5.91542053 C-3.24808548 5.01163162 -3.25030609 4.10784271 -3.25259399 3.17666626 C-3.08677921 0.34115132 -2.8362359 0.15995116 0 0 Z " fill="#EFEFEF" transform="translate(973.1323394775391,158.87974548339844)"/>
<path d="M0 0 C1.40897804 0.00333092 1.40897804 0.00333092 2.84642029 0.00672913 C3.90744461 0.00680466 4.96846893 0.00688019 6.06164551 0.00695801 C7.21579453 0.01211929 8.36994354 0.01728058 9.55906677 0.02259827 C10.73404221 0.02401321 11.90901764 0.02542816 13.11959839 0.02688599 C16.88981116 0.0325046 20.65996556 0.04506026 24.43016052 0.05775452 C26.97898779 0.06276712 29.52781599 0.06733044 32.0766449 0.07142639 C38.34035761 0.0816312 44.60394336 0.10120299 50.86766052 0.12025452 C50.86766052 17.28025452 50.86766052 34.44025452 50.86766052 52.12025452 C43.33791913 52.14315674 35.80829761 52.1630859 28.27854919 52.17518616 C25.71474296 52.18022822 23.15093961 52.18706166 20.58714294 52.19569397 C16.91111031 52.20776516 13.23511554 52.21348394 9.55906677 52.21791077 C8.40491776 52.22307205 7.25076874 52.22823334 6.06164551 52.23355103 C5.00062119 52.23362656 3.93959686 52.23370209 2.84642029 52.23377991 C1.90710159 52.23600052 0.9677829 52.23822113 0 52.24050903 C-2.13233948 52.12025452 -2.13233948 52.12025452 -3.13233948 51.12025452 C-3.23080914 49.56026404 -3.26032565 47.99584907 -3.26173401 46.43275452 C-3.26488617 45.43502014 -3.26803833 44.43728577 -3.27128601 43.40931702 C-3.26926178 42.32392639 -3.26723755 41.23853577 -3.26515198 40.12025452 C-3.2661087 39.01423889 -3.26706543 37.90822327 -3.26805115 36.76869202 C-3.26873314 34.42494144 -3.26687752 32.08118899 -3.26271057 29.73744202 C-3.25736262 26.13583664 -3.26265494 22.53435598 -3.26905823 18.93275452 C-3.26839745 16.66192091 -3.26711629 14.39108737 -3.26515198 12.12025452 C-3.26717621 11.03486389 -3.26920044 9.94947327 -3.27128601 8.83119202 C-3.26813385 7.83345764 -3.26498169 6.83572327 -3.26173401 5.80775452 C-3.26093842 4.9247467 -3.26014282 4.04173889 -3.25932312 3.13197327 C-3.08228729 0.32731047 -2.80658452 0.15827896 0 0 Z " fill="#EFF0EF" transform="translate(919.1323394775391,652.8797454833984)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.25394531 0.845625 1.50789063 1.69125 1.76953125 2.5625 C4.02209666 10.06445543 4.02209666 10.06445543 6.8125 17.375 C7.96931081 20.90631722 7.8530712 22.23508964 7.2644043 25.72998047 C6.66137976 30.90719387 6.94300272 36.17114816 7 41.375 C7.02536987 43.7369348 7.04645006 46.09892099 7.0625 48.4609375 C7.07410156 49.50040527 7.08570313 50.53987305 7.09765625 51.61083984 C7 54 7 54 6 55 C4.34261557 55.09346915 2.68125356 55.11744977 1.02124023 55.11352539 C-0.03978409 55.11344986 -1.10080841 55.11337433 -2.19398499 55.11329651 C-3.92520851 55.10555458 -3.92520851 55.10555458 -5.69140625 55.09765625 C-6.86638168 55.0962413 -8.04135712 55.09482635 -9.25193787 55.09336853 C-13.02215064 55.08774992 -16.79230504 55.07519426 -20.5625 55.0625 C-23.11132727 55.0574874 -25.66015547 55.05292408 -28.20898438 55.04882812 C-34.47269709 55.03862331 -40.73628284 55.01905152 -47 55 C-47 37.84 -47 20.68 -47 3 C-40.25 1.875 -40.25 1.875 -36.55517578 1.88647461 C-35.32457932 1.88658791 -35.32457932 1.88658791 -34.06912231 1.88670349 C-33.20326508 1.89186478 -32.33740784 1.89702606 -31.4453125 1.90234375 C-30.54376434 1.9037587 -29.64221619 1.90517365 -28.71334839 1.90663147 C-25.850531 1.9122026 -22.98779352 1.92474974 -20.125 1.9375 C-18.17708447 1.94251873 -16.2291677 1.94708099 -14.28125 1.95117188 C-9.52080282 1.96216258 -4.76041493 1.97940723 0 2 C0 1.34 0 0.68 0 0 Z " fill="#EFEFEF" transform="translate(264,545)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.16 53 34.32 53 52 C47.58428233 52.67696471 42.80465373 53.12801012 37.421875 53.1328125 C36.72918518 53.13376923 36.03649536 53.13472595 35.32281494 53.13571167 C33.86739002 53.13638697 32.41196197 53.13457844 30.95654297 53.13037109 C28.76913409 53.12504658 26.5819336 53.1303214 24.39453125 53.13671875 C22.96614539 53.13605722 21.53775966 53.13477451 20.109375 53.1328125 C18.20623535 53.13112061 18.20623535 53.13112061 16.26464844 53.12939453 C10.83254387 52.96457799 5.41583192 52.45131933 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFF0EF" transform="translate(810,653)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.16 53 34.32 53 52 C35.51 52 18.02 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFF0EF" transform="translate(917,865)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.16 53 34.32 53 52 C35.51 52 18.02 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#EFEFEF" transform="translate(863,706)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.16 53 34.32 53 52 C35.51 52 18.02 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#F0F0F0" transform="translate(702,653)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 17.16 53 34.32 53 52 C35.51 52 18.02 52 0 52 C0 34.84 0 17.68 0 0 Z " fill="#FEFEFE" transform="translate(702,159)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C56.2876071 6.57521419 56.12449325 18.17571336 53.90234375 25.11328125 C52.92371651 27.70741491 51.80988492 30.23584777 50.703125 32.77734375 C48.59530623 37.69917228 47.37068803 42.80473737 46.125 48 C45.91020996 48.89195068 45.69541992 49.78390137 45.47412109 50.70288086 C44.97501026 52.8000943 44.48632056 54.89978379 44 57 C42 55 42 55 40 52 C39.67 52.33 39.34 52.66 39 53 C36.20006403 53.10103255 33.42531356 53.13970088 30.625 53.1328125 C29.78533691 53.13376923 28.94567383 53.13472595 28.08056641 53.13571167 C26.30175705 53.13639348 24.52294523 53.13453917 22.74414062 53.13037109 C20.01166224 53.12502283 17.27934824 53.13031605 14.546875 53.13671875 C12.8229163 53.13605797 11.09895771 53.13477681 9.375 53.1328125 C8.55209473 53.13483673 7.72918945 53.13686096 6.88134766 53.13894653 C1.11495054 53.11495054 1.11495054 53.11495054 0 52 C-0.09340434 50.37325222 -0.11745171 48.74245949 -0.11352539 47.11303711 C-0.11340454 46.05741577 -0.11328369 45.00179443 -0.11315918 43.91418457 C-0.10548523 42.23769836 -0.10548523 42.23769836 -0.09765625 40.52734375 C-0.09664917 39.50612427 -0.09564209 38.48490479 -0.09460449 37.43273926 C-0.08935415 33.60098149 -0.07539303 29.76923967 -0.0625 25.9375 C-0.0315625 13.0984375 -0.0315625 13.0984375 0 0 Z " fill="#EFF0F0" transform="translate(217,369)"/>
<path d="M0 0 C0.81082031 -0.00257813 1.62164063 -0.00515625 2.45703125 -0.0078125 C5.71857101 0.15083178 8.9549231 0.6632033 12.1875 1.125 C12.1875 18.615 12.1875 36.105 12.1875 54.125 C-5.3025 54.125 -22.7925 54.125 -40.8125 54.125 C-41.8125 45.125 -41.8125 45.125 -40.3996582 42.81030273 C-39.70702881 42.25286377 -39.01439941 41.6954248 -38.30078125 41.12109375 C-33.83733302 37.19484959 -30.47181379 32.99624815 -27 28.1875 C-26.40396973 27.3742627 -25.80793945 26.56102539 -25.19384766 25.72314453 C-20.62803432 19.42794871 -16.36397837 12.96277218 -12.36401367 6.29321289 C-9.27118157 1.28303079 -9.27118157 1.28303079 -6.81420898 0.43652344 C-4.5146485 0.07864575 -2.32765372 -0.00733119 0 0 Z " fill="#FCFDFD" transform="translate(742.8125,598.875)"/>
<path d="M0 0 C-0.78375 1.03125 -1.5675 2.0625 -2.375 3.125 C-3.58637594 4.74773312 -4.79425115 6.37308139 -6 8 C-6.73863281 8.99515625 -7.47726562 9.9903125 -8.23828125 11.015625 C-18.1719118 24.56570216 -26.83827093 38.79660244 -34 54 C-36.97 53.34 -39.94 52.68 -43 52 C-43 34.84 -43 17.68 -43 0 C-37.204375 -0.185625 -31.40875 -0.37125 -25.4375 -0.5625 C-23.6217749 -0.62381104 -21.8060498 -0.68512207 -19.93530273 -0.74829102 C-18.47641411 -0.79230819 -17.01751182 -0.83587601 -15.55859375 -0.87890625 C-14.81710083 -0.90561401 -14.07560791 -0.93232178 -13.31164551 -0.95983887 C-8.73949496 -1.08774707 -4.51049907 -0.77211425 0 0 Z " fill="#EEEFEF" transform="translate(314,317)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C57.13404247 6.26808495 55 13.99206799 55 21 C36.85 21 18.7 21 0 21 C0 14.07 0 7.14 0 0 Z " fill="#EFEFEF" transform="translate(0,473)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53.33 12.87 53.66 25.74 54 39 C53.34 39 52.68 39 52 39 C52.495 40.98 52.495 40.98 53 43 C52.01 43.495 52.01 43.495 51 44 C50.66871094 43.58492188 50.33742188 43.16984375 49.99609375 42.7421875 C37.96127732 28.32453774 23.05233211 16.69507589 7.71142578 6.03466797 C7.00228027 5.54111816 6.29313477 5.04756836 5.5625 4.5390625 C4.92441406 4.09771973 4.28632812 3.65637695 3.62890625 3.20166016 C2 2 2 2 0 0 Z " fill="#EDEFEE" transform="translate(648,264)"/>
<path d="M0 0 C17.49 0 34.98 0 53 0 C53 4.29 53 8.58 53 13 C53.99 13.33 54.98 13.66 56 14 C55.08347656 14.14695313 55.08347656 14.14695313 54.1484375 14.296875 C50.76309107 14.84997385 47.38116889 15.42203551 44 16 C42.76950928 16.20931152 42.76950928 16.20931152 41.51416016 16.42285156 C30.89346494 18.24420508 20.47001246 20.25452306 10.09765625 23.18359375 C6.38214196 24.16284027 2.82360488 24.68786899 -1 25 C-1 24.34 -1 23.68 -1 23 C-2.32 23 -3.64 23 -5 23 C-5 22.34 -5 21.68 -5 21 C-3.68 20.67 -2.36 20.34 -1 20 C-0.67 13.4 -0.34 6.8 0 0 Z " fill="#FCFDFD" transform="translate(433,211)"/>
<path d="M0 0 C-0.96486328 0.58394531 -0.96486328 0.58394531 -1.94921875 1.1796875 C-19.24777166 11.88949059 -34.93061974 25.33474011 -49 40 C-50.32419476 35.99914344 -50.14384587 31.93204911 -50.1328125 27.76953125 C-50.13376923 26.9785051 -50.13472595 26.18747894 -50.13571167 25.3724823 C-50.13639066 23.70575887 -50.134556 22.03903277 -50.13037109 20.37231445 C-50.12499748 17.81130102 -50.13033648 15.25046127 -50.13671875 12.68945312 C-50.13605834 11.07031211 -50.13477794 9.45117121 -50.1328125 7.83203125 C-50.13483673 7.0622847 -50.13686096 6.29253815 -50.13894653 5.49946594 C-50.11496553 0.11496553 -50.11496553 0.11496553 -49 -1 C-47.5384677 -1.13268003 -46.07080256 -1.19877091 -44.60375977 -1.23706055 C-43.20209312 -1.27666145 -43.20209312 -1.27666145 -41.77210999 -1.31706238 C-40.75547775 -1.34004898 -39.73884552 -1.36303558 -38.69140625 -1.38671875 C-37.65435043 -1.41224319 -36.61729462 -1.43776764 -35.54881287 -1.46406555 C-33.35055485 -1.51617647 -31.15223155 -1.56559077 -28.95385742 -1.61254883 C-25.58020144 -1.68710879 -22.20722049 -1.77773236 -18.83398438 -1.86914062 C-16.70314727 -1.91765499 -14.57228814 -1.96521299 -12.44140625 -2.01171875 C-11.42679825 -2.04077805 -10.41219025 -2.06983734 -9.36683655 -2.09977722 C-8.42923996 -2.11672134 -7.49164337 -2.13366547 -6.52563477 -2.15112305 C-5.69814224 -2.17031296 -4.87064972 -2.18950287 -4.01808167 -2.20927429 C-2 -2 -2 -2 0 0 Z " fill="#EDF0F0" transform="translate(374,265)"/>
<path d="M0 0 C1.4540625 0.0309375 1.4540625 0.0309375 2.9375 0.0625 C4.29835719 2.78421438 4.16451682 5.15032141 4.3125 8.1875 C4.86459547 15.88286148 6.19927223 22.47527822 11.9375 28.0625 C18.92705134 32.61473547 25.50518512 35.37225305 33.9375 34.0625 C42.7819134 30.81880016 48.04558992 27.12334264 52.6875 19 C54.50579186 14.48982355 54.44649468 9.6589735 54.62890625 4.85546875 C54.9375 2.0625 54.9375 2.0625 56.9375 0.0625 C59.5625 -0.0625 59.5625 -0.0625 61.9375 0.0625 C64.50610043 5.19970087 63.48238708 12.6525423 62.25390625 18.0859375 C59.00227099 27.71941292 54.38054104 33.72329888 45.59765625 38.8359375 C36.59084468 42.98885796 26.03520607 43.89111653 16.51171875 41.03515625 C7.58591877 36.94085664 0.28486808 30.08684417 -3.44921875 20.875 C-4.85626899 14.42228551 -4.50889507 7.61938499 -4.0625 1.0625 C-3.0625 0.0625 -3.0625 0.0625 0 0 Z " fill="#FBF7F4" transform="translate(482.0625,488.9375)"/>
<path d="M0 0 C0 7.92 0 15.84 0 24 C-17.49 24 -34.98 24 -53 24 C-53 24.66 -53 25.32 -53 26 C-53.66 26 -54.32 26 -55 26 C-53.4943193 22.16735822 -51.23168738 20.462238 -48 18 C-47.44441406 17.37996094 -46.88882812 16.75992187 -46.31640625 16.12109375 C-43.2728321 13.33414474 -40.0380162 11.78291128 -36.3125 10.0625 C-35.57225586 9.71695068 -34.83201172 9.37140137 -34.06933594 9.01538086 C-23.56076862 4.26525137 -11.60133208 0 0 0 Z " fill="#F8FDFC" transform="translate(486,345)"/>
<path d="M0 0 C1.08809212 0.00212242 1.08809212 0.00212242 2.19816589 0.00428772 C4.50064325 0.00985694 6.8030211 0.02240364 9.10546875 0.03515625 C10.67252463 0.04017523 12.23958205 0.04473744 13.80664062 0.04882812 C17.63548526 0.05896271 21.46411644 0.07854384 25.29296875 0.09765625 C25.62296875 8.67765625 25.95296875 17.25765625 26.29296875 26.09765625 C25.96296875 26.09765625 25.63296875 26.09765625 25.29296875 26.09765625 C25.29296875 24.44765625 25.29296875 22.79765625 25.29296875 21.09765625 C12.75296875 21.09765625 0.21296875 21.09765625 -12.70703125 21.09765625 C-12.70703125 14.49765625 -12.70703125 7.89765625 -12.70703125 1.09765625 C-8.32747449 0.2217449 -4.41742737 -0.03275672 0 0 Z " fill="#EFEFEF" transform="translate(229.70703125,472.90234375)"/>
<path d="M0 0 C11.55 0 23.1 0 35 0 C34.67 5.61 34.34 11.22 34 17 C33.9628207 20.13700358 33.93834817 23.24308712 34 26.375 C34.13146552 33.60560345 34.13146552 33.60560345 33 37 C19.28219864 30.56978061 6.1101768 16.31960344 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#FCFBFB" transform="translate(399,547)"/>
<path d="M0 0 C17.82 0 35.64 0 54 0 C54 4.95 54 9.9 54 15 C46.79163272 14.8818923 39.58340735 14.75765377 32.37524414 14.62768555 C29.92214851 14.58432398 27.46902247 14.54264981 25.01586914 14.50268555 C21.49355899 14.44501279 17.97140216 14.38130948 14.44921875 14.31640625 C13.34913986 14.29969376 12.24906097 14.28298126 11.11564636 14.26576233 C9.58439873 14.2358445 9.58439873 14.2358445 8.0222168 14.20532227 C7.12286911 14.18977798 6.22352142 14.1742337 5.29692078 14.15821838 C3 14 3 14 0 13 C0 8.71 0 4.42 0 0 Z " fill="#EBEDED" transform="translate(486,211)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C0.67 15.84 0.34 31.68 0 48 C-6.93 48 -13.86 48 -21 48 C-19.845 45.751875 -18.69 43.50375 -17.5 41.1875 C-10.76775746 27.85685118 -5.22144298 13.98242183 0 0 Z " fill="#EAEEED" transform="translate(755,552)"/>
<path d="M0 0 C23.47027881 4.51459365 48.46257366 12.91018651 68 27 C67.34 27.33 66.68 27.66 66 28 C63.64018187 27.06421005 61.30368736 26.06652192 59 25 C59 24.34 59 23.68 59 23 C58.31292969 23.02320313 57.62585938 23.04640625 56.91796875 23.0703125 C55.56638672 23.09738281 55.56638672 23.09738281 54.1875 23.125 C53.29417969 23.14820313 52.40085937 23.17140625 51.48046875 23.1953125 C49 23 49 23 46 21 C46.66 20.34 47.32 19.68 48 19 C45.525 18.01 45.525 18.01 43 17 C43 16.34 43 15.68 43 15 C42.32453125 15.02320313 41.6490625 15.04640625 40.953125 15.0703125 C39.61507812 15.09738281 39.61507812 15.09738281 38.25 15.125 C36.92742188 15.15980469 36.92742188 15.15980469 35.578125 15.1953125 C32.8864142 14.99139502 31.30095026 14.36551721 29 13 C29.99 13 30.98 13 32 13 C32 12.34 32 11.68 32 11 C31.39671875 10.87882812 30.7934375 10.75765625 30.171875 10.6328125 C29.37265625 10.46523438 28.5734375 10.29765625 27.75 10.125 C26.96109375 9.96257812 26.1721875 9.80015625 25.359375 9.6328125 C23 9 23 9 21.03125 7.9375 C18.47659974 6.75843065 16.5488555 6.80134591 13.75 6.875 C12.41195312 6.90207031 12.41195312 6.90207031 11.046875 6.9296875 C10.37140625 6.95289063 9.6959375 6.97609375 9 7 C8.67 6.34 8.34 5.68 8 5 C8.33 4.34 8.66 3.68 9 3 C8.2575 3.37125 7.515 3.7425 6.75 4.125 C4 5 4 5 1.6875 4.125 C1.130625 3.75375 0.57375 3.3825 0 3 C0 2.01 0 1.02 0 0 Z " fill="#D14674" transform="translate(553,265)"/>
<path d="M0 0 C3.45826342 -0.05789006 6.91640293 -0.09355821 10.375 -0.125 C11.35984375 -0.14175781 12.3446875 -0.15851563 13.359375 -0.17578125 C14.77089844 -0.18544922 14.77089844 -0.18544922 16.2109375 -0.1953125 C17.08024902 -0.20578613 17.94956055 -0.21625977 18.84521484 -0.22705078 C21 0 21 0 23 2 C23.5 4.1875 23.5 4.1875 23 7 C21.25247516 9.58376373 19.32164007 11.91292979 17 14 C16.34 14 15.68 14 15 14 C15 14.66 15 15.32 15 16 C13.7421875 17.23657227 13.7421875 17.23657227 11.875 18.75390625 C5.2090302 24.42203798 -0.83897236 30.73363132 -7 36.9375 C-8.2640885 38.20661373 -9.52840956 39.47549589 -10.79296875 40.74414062 C-13.86466724 43.8267632 -16.93320008 46.91250428 -20 50 C-20.495 48.515 -20.495 48.515 -21 47 C-19.71034824 45.62437146 -18.37310707 44.29233607 -17 43 C-16.34 43 -15.68 43 -15 43 C-15 42.34 -15 41.68 -15 41 C-14.34 41 -13.68 41 -13 41 C-13 40.34 -13 39.68 -13 39 C-12.34 39 -11.68 39 -11 39 C-11 38.34 -11 37.68 -11 37 C-10.34 37 -9.68 37 -9 37 C-9 36.34 -9 35.68 -9 35 C-8.34 35 -7.68 35 -7 35 C-6.896875 34.360625 -6.79375 33.72125 -6.6875 33.0625 C-6.460625 32.381875 -6.23375 31.70125 -6 31 C-5.01 30.67 -4.02 30.34 -3 30 C-3 29.34 -3 28.68 -3 28 C-1.29059971 26.39771617 0.53301528 24.98705258 2.37109375 23.53515625 C4.26558258 21.99243114 4.26558258 21.99243114 5 19 C5.99 18.67 6.98 18.34 8 18 C9.00642948 16.67151309 10.00692179 15.33849671 11 14 C11.66 14 12.32 14 13 14 C13.33 13.01 13.66 12.02 14 11 C14.99 11 15.98 11 17 11 C17 10.34 17 9.68 17 9 C17.66 9 18.32 9 19 9 C19.6814823 7.10820797 19.6814823 7.10820797 20 5 C16.38260457 1.38260457 12.74358778 1.69396274 7.875 1.4375 C7.12089844 1.39431641 6.36679687 1.35113281 5.58984375 1.30664062 C3.72678112 1.2005168 1.86341476 1.09974999 0 1 C0 0.67 0 0.34 0 0 Z " fill="#D74F7D" transform="translate(720,446)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.15410894 8.76237448 1.30228743 17.52482359 1.4429636 26.28742409 C1.50847488 30.35654809 1.57600353 34.42561747 1.64819336 38.49462891 C1.71782723 42.42380453 1.78209548 46.3530351 1.84269524 50.28236008 C1.86671091 51.77903791 1.89263705 53.27568639 1.92053413 54.77229691 C1.95937352 56.87370469 1.99132631 58.97511565 2.02172852 61.07666016 C2.04171402 62.27134918 2.06169952 63.46603821 2.08229065 64.69692993 C2.00259131 67.89598725 1.60937149 70.86261045 1 74 C0.67 74 0.34 74 0 74 C0 72.02 0 70.04 0 68 C-17.16 68 -34.32 68 -52 68 C-52 67.67 -52 67.34 -52 67 C-34.84 67 -17.68 67 0 67 C0 49.84 0 32.68 0 15 C-6.6 15 -13.2 15 -20 15 C-20 14.67 -20 14.34 -20 14 C-13.4 14 -6.8 14 0 14 C0 9.38 0 4.76 0 0 Z " fill="#F6F6F6" transform="translate(162,480)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C2 0.66 2 1.32 2 2 C2.66 2 3.32 2 4 2 C4.33 2.66 4.66 3.32 5 4 C5.99 3.67 6.98 3.34 8 3 C8.33 4.65 8.66 6.3 9 8 C11.31 8.66 13.62 9.32 16 10 C15.95875 10.78375 15.9175 11.5675 15.875 12.375 C15.71271266 15.16116119 15.71271266 15.16116119 18 17 C19.98821313 17.39764263 21.98944339 17.73775349 24 18 C24.061875 18.94875 24.12375 19.8975 24.1875 20.875 C24.455625 21.90625 24.72375 22.9375 25 24 C27.47590076 25.39666197 29.16264185 26 32 26 C32.66 28.31 33.32 30.62 34 33 C35.98 33 37.96 33 40 33 C40 35.31 40 37.62 40 40 C36.83199926 38.59779351 34.68824332 36.94085834 32.24121094 34.5 C31.52076599 33.78585937 30.80032104 33.07171875 30.05804443 32.3359375 C28.90782806 31.17964844 28.90782806 31.17964844 27.734375 30 C26.94097717 29.20851563 26.14757935 28.41703125 25.33013916 27.6015625 C23.65675946 25.92954263 21.98589819 24.25499903 20.31738281 22.578125 C17.75286403 20.00287602 15.17783011 17.43848948 12.6015625 14.875 C10.97852473 13.25064116 9.35610719 11.62566231 7.734375 10 C6.95946716 9.22914063 6.18455933 8.45828125 5.38616943 7.6640625 C4.67833313 6.94992187 3.97049683 6.23578125 3.24121094 5.5 C2.61373962 4.8709375 1.98626831 4.241875 1.33978271 3.59375 C0 2 0 2 0 0 Z " fill="#A12760" transform="translate(616,454)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1 2.64 1 5.28 1 8 C10.9 8 20.8 8 31 8 C31 8.33 31 8.66 31 9 C21.1 9 11.2 9 1 9 C1.08378906 12.22265625 1.16757813 15.4453125 1.25390625 18.765625 C2.02562196 50.54485235 1.86998459 82.22484837 1 114 C0.67 114 0.34 114 0 114 C-0.15401963 100.31754627 -0.30219936 86.63504288 -0.4429636 72.95244598 C-0.50851154 66.598796 -0.5760563 60.24518042 -0.64819336 53.89160156 C-0.71776025 47.75788103 -0.78204416 41.62412562 -0.84269524 35.49031067 C-0.86673529 33.15238949 -0.89266558 30.81448695 -0.92053413 28.47660828 C-0.95929895 25.19732575 -0.99128865 21.91804081 -1.02172852 18.63867188 C-1.03467453 17.6762558 -1.04762054 16.71383972 -1.06095886 15.72225952 C-1.10263324 10.37702915 -0.79068443 5.28835992 0 0 Z " fill="#F6F7F6" transform="translate(162,697)"/>
<path d="M0 0 C1.91914553 0.93241504 3.83522386 1.87114475 5.75 2.8125 C6.81734375 3.33457031 7.8846875 3.85664063 8.984375 4.39453125 C11.55233242 5.7616692 13.74470783 7.17715463 16 9 C15.67 9.99 15.34 10.98 15 12 C13.67696283 12.3721042 12.34262065 12.70630173 11 13 C10.67 13.66 10.34 14.32 10 15 C5.22390502 13.35821735 1.20617096 10.73453298 -3 8 C-2.5359375 7.13375 -2.5359375 7.13375 -2.0625 6.25 C-1.07416636 4.15705816 -0.4831387 2.25464725 0 0 Z " fill="#DCE0DF" transform="translate(630,266)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C2.48572053 11.51433409 3.19368943 22.88554126 3.1875 34.5 C3.18814453 35.65532227 3.18878906 36.81064453 3.18945312 38.00097656 C3.14291981 45.37650665 2.72411778 52.66049547 2 60 C1.67 60 1.34 60 1 60 C-0.05476516 54.83931509 -0.12969365 49.90287993 -0.09765625 44.6640625 C-0.0962413 43.78471039 -0.09482635 42.90535828 -0.09336853 41.99935913 C-0.08779877 39.20787058 -0.0752519 36.41646406 -0.0625 33.625 C-0.05748109 31.72526158 -0.05291887 29.8255219 -0.04882812 27.92578125 C-0.03783925 23.28382286 -0.02059557 18.64192531 0 14 C-0.33 14 -0.66 14 -1 14 C-0.67 9.38 -0.34 4.76 0 0 Z " fill="#2E6865" transform="translate(764,441)"/>
<path d="M0 0 C4.91734018 1.76282007 7.97009753 5.25126968 11.3125 9.1875 C11.3125 9.5175 11.3125 9.8475 11.3125 10.1875 C5.7025 10.1875 0.0925 10.1875 -5.6875 10.1875 C-5.6875 3.1875 -5.6875 3.1875 -4.5625 1.1875 C-2.6875 0.1875 -2.6875 0.1875 0 0 Z " fill="#9BDDC6" transform="translate(489.6875,248.8125)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.06058594 0.68964844 1.12117188 1.37929688 1.18359375 2.08984375 C1.26738281 3.02957031 1.35117187 3.96929687 1.4375 4.9375 C1.52644531 5.95328125 1.61539062 6.9690625 1.70703125 8.015625 C1.87614818 9.7383628 2.06864329 11.45982733 2.32421875 13.171875 C3.75358602 22.75049202 2.80853554 33.52327379 1 43 C0.01 43.495 0.01 43.495 -1 44 C-1.02491316 39.18026089 -1.04295998 34.36056015 -1.05493164 29.54077148 C-1.05992803 27.90469712 -1.06672739 26.26862715 -1.07543945 24.63256836 C-1.16225376 7.89783459 -1.16225376 7.89783459 0 0 Z " fill="#D2DCDB" transform="translate(267,445)"/>
<path d="M0 0 C0.99 0.495 0.99 0.495 2 1 C2 3.31 2 5.62 2 8 C2.66 7.01 3.32 6.02 4 5 C4.33 6.65 4.66 8.3 5 10 C5.33 10 5.66 10 6 10 C6 16.6 6 23.2 6 30 C5.01 30.33 4.02 30.66 3 31 C-0.58165209 9.39260417 -0.58165209 9.39260417 0 0 Z " fill="#DCE2E2" transform="translate(266,490)"/>
<path d="M0 0 C0 0.66 0 1.32 0 2 C-1.28463135 2.42297363 -1.28463135 2.42297363 -2.59521484 2.85449219 C-5.82033779 3.91806413 -9.0444931 4.98447904 -12.26806641 6.05273438 C-13.65441681 6.51153122 -15.04112665 6.96924359 -16.42822266 7.42578125 C-24.38588327 10.04577637 -32.27400477 12.74379813 -40 16 C-39.67 15.01 -39.34 14.02 -39 13 C-37.02 12.67 -35.04 12.34 -33 12 C-32.67 11.01 -32.34 10.02 -32 9 C-31.34 8.9175 -30.68 8.835 -30 8.75 C-26.7101066 7.92752665 -24.10849827 6.6019765 -21.11328125 5.05078125 C-14.29611273 1.66109857 -7.67299752 -0.2256764 0 0 Z " fill="#E4F9F5" transform="translate(450,274)"/>
<path d="M0 0 C-3.00663043 2.00442028 -4.6438078 2.50017063 -8.125 3.125 C-9.45917969 3.37636719 -9.45917969 3.37636719 -10.8203125 3.6328125 C-14.89332927 4.10316087 -18.9052408 4.07147959 -23 4 C-22.97643433 4.88522339 -22.97643433 4.88522339 -22.95239258 5.78833008 C-22.89002061 8.46295586 -22.85100343 11.13742864 -22.8125 13.8125 C-22.77479492 15.2056543 -22.77479492 15.2056543 -22.73632812 16.62695312 C-22.72182617 17.9659668 -22.72182617 17.9659668 -22.70703125 19.33203125 C-22.68346558 20.56530151 -22.68346558 20.56530151 -22.65942383 21.82348633 C-23 24 -23 24 -24.3503418 25.8112793 C-26 27 -26 27 -28.6875 26.6875 C-29.450625 26.460625 -30.21375 26.23375 -31 26 C-29 23 -29 23 -26 22 C-24.88176185 19.76352369 -24.80603939 18.35108471 -24.68359375 15.8671875 C-24.64169922 15.06152344 -24.59980469 14.25585938 -24.55664062 13.42578125 C-24.51732422 12.58402344 -24.47800781 11.74226562 -24.4375 10.875 C-24.37272461 9.60076172 -24.37272461 9.60076172 -24.30664062 8.30078125 C-24.20045764 6.20071777 -24.09971503 4.10038052 -24 2 C-15.95072024 0.70098079 -8.16240568 -0.33853295 0 0 Z " fill="#D07296" transform="translate(561,679)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C3.31 3 5.62 3 8 3 C9.35306884 7.05920652 7.84599602 9.41865449 6.1875 13.125 C5.91357422 13.77082031 5.63964844 14.41664063 5.35742188 15.08203125 C3.26584507 19.86707746 3.26584507 19.86707746 1 21 C0.67 14.07 0.34 7.14 0 0 Z " fill="#F5F8F8" transform="translate(270,366)"/>
<path d="M0 0 C0.66 0.66 1.32 1.32 2 2 C1.5399605 5.9521575 0.26252789 9.75751331 -0.875 13.5625 C-1.20242188 14.67753906 -1.52984375 15.79257812 -1.8671875 16.94140625 C-2.92484384 19.79707836 -4.03488285 21.70362025 -6 24 C-5.34 24.33 -4.68 24.66 -4 25 C-7 29.5 -7 29.5 -10 34 C-8.46680366 22.02573659 -4.98126903 10.96287487 0 0 Z " fill="#35C3A2" transform="translate(303,406)"/>
<path d="M0 0 C0.86803253 0.35190651 0.86803253 0.35190651 1.75360107 0.71092224 C0.70172607 1.23685974 0.70172607 1.23685974 -0.37139893 1.77342224 C-3.49392587 3.87773387 -5.41804197 6.13668856 -7.78155518 9.02342224 C-9.24639893 10.71092224 -9.24639893 10.71092224 -11.68389893 12.64842224 C-13.98478155 14.50035216 -15.66131591 16.28238528 -17.55889893 18.52342224 C-20.60022679 22.09598642 -23.88945644 25.09158629 -27.46514893 28.11717224 C-29.68545977 30.10376616 -31.41183121 32.37026688 -33.24639893 34.71092224 C-34.87996843 36.08460569 -36.53889913 37.43029739 -38.24639893 38.71092224 C-38.90639893 38.38092224 -39.56639893 38.05092224 -40.24639893 37.71092224 C-34.92537391 32.26343829 -29.58508985 26.8354038 -24.23077393 21.42063904 C-22.41048821 19.57516186 -20.59470895 17.72522868 -18.7835083 15.87083435 C-16.1838236 13.2107084 -13.56851273 10.56687091 -10.94952393 7.92576599 C-10.13896545 7.08940109 -9.32840698 6.25303619 -8.49328613 5.3913269 C-7.73279968 4.6304628 -6.97231323 3.86959869 -6.18878174 3.0856781 C-5.52259827 2.40839157 -4.85641479 1.73110504 -4.17004395 1.03329468 C-2.24639893 -0.28907776 -2.24639893 -0.28907776 0 0 Z " fill="#EAF9F6" transform="translate(539.2463989257813,329.28907775878906)"/>
<path d="M0 0 C1.47919922 0.06960938 1.47919922 0.06960938 2.98828125 0.140625 C3.98214844 0.17671875 4.97601562 0.2128125 6 0.25 C7.13888672 0.31960938 7.13888672 0.31960938 8.30078125 0.390625 C4.09718033 3.70643494 -0.43848087 5.80943021 -5.26171875 8.078125 C-6.12474609 8.49384766 -6.98777344 8.90957031 -7.87695312 9.33789062 C-8.70646484 9.73041016 -9.53597656 10.12292969 -10.390625 10.52734375 C-11.14545166 10.88530029 -11.90027832 11.24325684 -12.67797852 11.61206055 C-14.69921875 12.390625 -14.69921875 12.390625 -17.69921875 12.390625 C-17.36921875 10.740625 -17.03921875 9.090625 -16.69921875 7.390625 C-15.93996094 7.22046875 -15.18070313 7.0503125 -14.3984375 6.875 C-12.90763672 6.51148438 -12.90763672 6.51148438 -11.38671875 6.140625 C-10.40058594 5.90859375 -9.41445313 5.6765625 -8.3984375 5.4375 C-5.58000958 4.62764839 -5.58000958 4.62764839 -4.19921875 2.296875 C-2.69921875 0.390625 -2.69921875 0.390625 0 0 Z " fill="#D8779B" transform="translate(613.69921875,657.609375)"/>
<path d="M0 0 C0.68513672 -0.00386719 1.37027344 -0.00773437 2.07617188 -0.01171875 C7.1841133 -0.00169335 7.1841133 -0.00169335 9.4375 1.125 C9.4375 1.785 9.4375 2.445 9.4375 3.125 C10.4275 3.455 11.4175 3.785 12.4375 4.125 C3.5275 4.125 -5.3825 4.125 -14.5625 4.125 C-9.42966353 0.27537264 -6.16514138 -0.03499607 0 0 Z " fill="#EEF9F8" transform="translate(351.5625,416.875)"/>
<path d="M0 0 C2.69473638 8.08420915 0.37904963 14.66873519 -2.8125 22.125 C-3.16892578 22.99253906 -3.52535156 23.86007812 -3.89257812 24.75390625 C-5.76284109 29.26312741 -7.74903495 33.66848996 -10 38 C-11.48356761 34.14272421 -10.31383511 31.78693649 -9 28 C-8.83142517 25.24934768 -8.83142517 25.24934768 -9 23 C-8.01 23 -7.02 23 -6 23 C-3.60061221 16.5652782 -2.32807977 10.4338677 -1.4296875 3.625 C-1 1 -1 1 0 0 Z " fill="#D46F96" transform="translate(722,528)"/>
<path d="M0 0 C4 0 4 0 5.9375 1.8125 C6.618125 2.534375 7.29875 3.25625 8 4 C8.9075 4.53625 9.815 5.0725 10.75 5.625 C11.4925 6.07875 12.235 6.5325 13 7 C13 7.66 13 8.32 13 9 C13.66 9 14.32 9 15 9 C14.95875 9.94875 14.9175 10.8975 14.875 11.875 C14.65026182 15.10244856 14.65026182 15.10244856 17 17 C16.67 17.99 16.34 18.98 16 20 C15.26394531 19.11957031 14.52789063 18.23914063 13.76953125 17.33203125 C12.78397631 16.15875156 11.79829234 14.98558023 10.8125 13.8125 C10.32974609 13.23435547 9.84699219 12.65621094 9.34960938 12.06054688 C7.04130899 9.31847192 4.72297028 6.68329738 2.13671875 4.19921875 C0 2 0 2 0 0 Z " fill="#B13566" transform="translate(553,279)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1 3.3 1 6.6 1 10 C6.61 10 12.22 10 18 10 C16.53787551 12.92424897 14.22537218 13.34147999 11.27734375 14.40234375 C7.76495361 15.32412024 4.61542291 15.19368337 1 15 C0.87625 14.360625 0.7525 13.72125 0.625 13.0625 C0.41875 12.381875 0.2125 11.70125 0 11 C-0.66 10.67 -1.32 10.34 -2 10 C-1.34 10 -0.68 10 0 10 C0 6.7 0 3.4 0 0 Z " fill="#F8F5F6" transform="translate(540,590)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.69918305 2.58067563 2.38461049 5.16372847 3.0625 7.75 C3.26166016 8.47960937 3.46082031 9.20921875 3.66601562 9.9609375 C5.33219296 16.39179738 5.33219296 16.39179738 4 20 C1.9375 21.25 1.9375 21.25 0 22 C-1.28923485 18.13229545 -1.14505706 14.46562684 -1.125 10.4375 C-1.12886719 9.65697266 -1.13273438 8.87644531 -1.13671875 8.07226562 C-1.12667749 2.25335498 -1.12667749 2.25335498 0 0 Z " fill="#D64674" transform="translate(713,410)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C-0.5436892 4.9913131 -4.73605498 7.50654225 -9.25 10.25 C-9.99507812 10.70890625 -10.74015625 11.1678125 -11.5078125 11.640625 C-13.33550829 12.76536087 -15.16734673 13.8833601 -17 15 C-17.33 13.68 -17.66 12.36 -18 11 C-14.52740334 7.96147792 -11.05694957 5.91367946 -6.92578125 3.953125 C-4.80123511 2.94663382 -4.80123511 2.94663382 -2.1875 1.1875 C-1.465625 0.795625 -0.74375 0.40375 0 0 Z " fill="#D7769A" transform="translate(641,643)"/>
<path d="M0 0 C2.31 0 4.62 0 7 0 C7.33 2.31 7.66 4.62 8 7 C10.31 7.33 12.62 7.66 15 8 C15.33 8.99 15.66 9.98 16 11 C16.65129797 12.34090759 17.31513275 13.67592331 18 15 C12.01424571 14.70340857 9.5210457 12.20385229 5.625 8.0625 C5.07972656 7.51142578 4.53445313 6.96035156 3.97265625 6.39257812 C0 2.29546523 0 2.29546523 0 0 Z " fill="#A42D62" transform="translate(658,496)"/>
<path d="M0 0 C-0.33 0.99 -0.66 1.98 -1 3 C-2.77734375 3.73046875 -2.77734375 3.73046875 -4.9375 4.1875 C-5.64777344 4.34605469 -6.35804688 4.50460937 -7.08984375 4.66796875 C-9 5 -9 5 -11 5 C-12.69156537 5.72969487 -14.38269162 6.46044695 -16.0703125 7.19921875 C-21.085622 9.28047067 -25.57635166 10.26456821 -31 10 C-27.47352579 6.47352579 -22.39578191 5.48424881 -17.75 3.875 C-16.71230469 3.50246094 -15.67460937 3.12992187 -14.60546875 2.74609375 C-13.09146484 2.21822266 -13.09146484 2.21822266 -11.546875 1.6796875 C-10.62745117 1.35726074 -9.70802734 1.03483398 -8.76074219 0.70263672 C-5.74459948 -0.06500201 -3.09976736 -0.12264446 0 0 Z " fill="#4BC69D" transform="translate(449,277)"/>
<path d="M0 0 C2.29370117 0.42578125 2.29370117 0.42578125 4.29370117 2.42578125 C4.41870117 5.55078125 4.41870117 5.55078125 4.29370117 8.42578125 C3.63370117 7.10578125 2.97370117 5.78578125 2.29370117 4.42578125 C-7.86459597 4.67973868 -15.99104358 16.59942803 -22.70629883 23.42578125 C-23.36629883 23.09578125 -24.02629883 22.76578125 -24.70629883 22.42578125 C-21.6808368 19.27659012 -18.6391764 16.14425668 -15.58154297 13.02636719 C-14.54407273 11.96377464 -13.511137 10.89673484 -12.48291016 9.82519531 C-11.00271899 8.28425269 -9.50687266 6.76012246 -8.00708008 5.23828125 C-7.11158447 4.31660156 -6.21608887 3.39492188 -5.29345703 2.4453125 C-2.70629883 0.42578125 -2.70629883 0.42578125 0 0 Z " fill="#A13167" transform="translate(530.706298828125,579.57421875)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C3.125 6.75 3.125 6.75 2 9 C4.97 9.495 4.97 9.495 8 10 C8 10.99 8 11.98 8 13 C3.14036821 12.39254603 -0.7405518 10.27241033 -5 8 C-3.8141763 4.62496331 -2.72426311 2.35277269 0 0 Z " fill="#A52D68" transform="translate(565,343)"/>
<path d="M0 0 C4.92127034 -0.16682272 8.50343896 -0.24828052 13 2 C10.39902318 3.30048841 7.86044938 3.56471422 5 4 C5.66 5.65 6.32 7.3 7 9 C7.99 9 8.98 9 10 9 C10 9.66 10 10.32 10 11 C10.66 11 11.32 11 12 11 C13.625 13.5 13.625 13.5 15 16 C12 16 12 16 10.55786133 14.85424805 C10.0708374 14.32871338 9.58381348 13.80317871 9.08203125 13.26171875 C8.55029297 12.68873047 8.01855469 12.11574219 7.47070312 11.52539062 C6.92349609 10.91888672 6.37628906 10.31238281 5.8125 9.6875 C5.25369141 9.09259766 4.69488281 8.49769531 4.11914062 7.88476562 C0 3.38338484 0 3.38338484 0 0 Z " fill="#C8416B" transform="translate(539,263)"/>
<path d="M0 0 C5.93148406 5.65772326 10.65304739 12.51857651 14 20 C13.01 20.33 12.02 20.66 11 21 C8 16.25 8 16.25 8 14 C7.01 13.67 6.02 13.34 5 13 C4.690625 12.21625 4.38125 11.4325 4.0625 10.625 C2.85791386 7.64896365 1.66841391 6.68999547 -1 5 C-0.67 3.35 -0.34 1.7 0 0 Z " fill="#D2DFDD" transform="translate(705,330)"/>
<path d="M0 0 C3.45826342 -0.05789006 6.91640293 -0.09355821 10.375 -0.125 C11.35984375 -0.14175781 12.3446875 -0.15851563 13.359375 -0.17578125 C14.77089844 -0.18544922 14.77089844 -0.18544922 16.2109375 -0.1953125 C17.51490479 -0.21102295 17.51490479 -0.21102295 18.84521484 -0.22705078 C21 0 21 0 23 2 C23.5 4.1875 23.5 4.1875 23 7 C21.25247516 9.58376373 19.32164007 11.91292979 17 14 C16.34 14 15.68 14 15 14 C14.67 14.66 14.34 15.32 14 16 C14.61277612 13.03824877 15.25372522 11.61941217 17 9 C17.66 9 18.32 9 19 9 C19.6814823 7.10820797 19.6814823 7.10820797 20 5 C16.38260457 1.38260457 12.74358778 1.69396274 7.875 1.4375 C7.12089844 1.39431641 6.36679687 1.35113281 5.58984375 1.30664062 C3.72678112 1.2005168 1.86341476 1.09974999 0 1 C0 0.67 0 0.34 0 0 Z " fill="#DA678D" transform="translate(720,446)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.625 2.8125 1.625 2.8125 2 6 C1.34 6.99 0.68 7.98 0 9 C0 8.01 0 7.02 0 6 C-18.15 6 -36.3 6 -55 6 C-55 5.67 -55 5.34 -55 5 C-36.85 5 -18.7 5 0 5 C0 3.35 0 1.7 0 0 Z " fill="#F6F6F5" transform="translate(809,364)"/>
<path d="M0 0 C1 2 1 2 0.3125 4.5625 C-1 7 -1 7 -3.125 7.8125 C-3.74375 7.874375 -4.3625 7.93625 -5 8 C-5 8.66 -5 9.32 -5 10 C-5.99 10.66 -6.98 11.32 -8 12 C-8.73606499 15.56769552 -8.73606499 15.56769552 -9 19 C-10.65 18.67 -12.3 18.34 -14 18 C-13.75898603 12.43572085 -10.23981113 9.78146531 -6.4375 6.1875 C-5.82197266 5.59001953 -5.20644531 4.99253906 -4.57226562 4.37695312 C-3.05706751 2.9087379 -1.52969562 1.45310447 0 0 Z " fill="#9A2D67" transform="translate(489,619)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C1 3 1 3 -1 4 C-1.65213292 6.02463255 -1.65213292 6.02463255 -2 8 C-8.625 9 -8.625 9 -12 9 C-12.66 9.66 -13.32 10.32 -14 11 C-15.32 10.34 -16.64 9.68 -18 9 C-12 6 -6 3 0 0 Z " fill="#DCE2E1" transform="translate(410,256)"/>
<path d="M0 0 C1.95273962 2.92910944 2.75396363 5.08132291 3.6875 8.4375 C3.95949219 9.38496094 4.23148438 10.33242188 4.51171875 11.30859375 C5.00264436 14.01457569 5.03759439 15.47442685 4 18 C1.9375 19.25 1.9375 19.25 0 20 C-1.87457064 13.40924767 -1.13537936 6.67035373 0 0 Z M0 11 C0 12.65 0 14.3 0 16 C0.33 16 0.66 16 1 16 C1 14.35 1 12.7 1 11 C0.67 11 0.34 11 0 11 Z " fill="#D2DEDB" transform="translate(745,405)"/>
<path d="M0 0 C-1 1 -1 1 -2.85766602 1.11352539 C-3.64842529 1.10828857 -4.43918457 1.10305176 -5.25390625 1.09765625 C-6.10791016 1.09443359 -6.96191406 1.09121094 -7.84179688 1.08789062 C-8.73962891 1.07951172 -9.63746094 1.07113281 -10.5625 1.0625 C-11.46419922 1.05798828 -12.36589844 1.05347656 -13.29492188 1.04882812 C-15.53001314 1.03700225 -17.76497437 1.0205222 -20 1 C-20 0.01 -20 -0.98 -20 -2 C-13.2641942 -3.31787505 -5.88621186 -3.92414124 0 0 Z " fill="#F6F8F8" transform="translate(467,727)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C-0.32346506 5.0065438 -1.65729179 7.00628175 -3 9 C-3 10.32 -3 11.64 -3 13 C-3.66 13 -4.32 13 -5 13 C-5.10183594 13.58265625 -5.20367187 14.1653125 -5.30859375 14.765625 C-6.11517153 17.37219275 -7.24157009 18.73535414 -9.0625 20.75 C-9.61035156 21.36359375 -10.15820312 21.9771875 -10.72265625 22.609375 C-11.14417969 23.06828125 -11.56570313 23.5271875 -12 24 C-12.33 23.34 -12.66 22.68 -13 22 C-11.67948953 19.34109405 -10.30556706 16.80954352 -8.8125 14.25 C-8.41224609 13.54617188 -8.01199219 12.84234375 -7.59960938 12.1171875 C-5.21830427 7.96437665 -2.70234735 3.95101819 0 0 Z " fill="#CFDBDA" transform="translate(304,348)"/>
<path d="M0 0 C1.32 0.33 2.64 0.66 4 1 C2.59902171 3.65527296 1.18061525 6.29826152 -0.25 8.9375 C-0.64574219 9.69224609 -1.04148437 10.44699219 -1.44921875 11.22460938 C-1.84238281 11.94326172 -2.23554687 12.66191406 -2.640625 13.40234375 C-2.99672852 14.06741943 -3.35283203 14.73249512 -3.71972656 15.41772461 C-5.3253581 17.40210638 -6.52169666 17.63191251 -9 18 C-8.52354792 13.71193127 -7.34097516 11.73352513 -4 9 C-3.34 9 -2.68 9 -2 9 C-2.04125 8.071875 -2.0825 7.14375 -2.125 6.1875 C-2 3 -2 3 0 0 Z " fill="#D2DCD8" transform="translate(724,589)"/>
<path d="M0 0 C1.94566951 3.47547073 2.07637127 5.12506344 1 9 C0.34 9 -0.32 9 -1 9 C-1.2475 9.99 -1.495 10.98 -1.75 12 C-2.95812141 16.28095196 -4.90821294 20.09059215 -7 24 C-7.66 24 -8.32 24 -9 24 C-6.80148049 15.63019764 -3.50929804 7.88172441 0 0 Z " fill="#C7D6D5" transform="translate(287,378)"/>
<path d="M0 0 C-0.75 1.9375 -0.75 1.9375 -2 4 C-5.75515022 5.5887174 -9.33064022 4.67943626 -13.25 4.0625 C-14.51328125 3.86785156 -15.7765625 3.67320312 -17.078125 3.47265625 C-18.04234375 3.31667969 -19.0065625 3.16070313 -20 3 C-20 2.67 -20 2.34 -20 2 C-17.41842632 1.46867611 -14.83538244 0.94965621 -12.25 0.4375 C-11.52039063 0.28603516 -10.79078125 0.13457031 -10.0390625 -0.02148438 C-6.33442927 -0.74557178 -3.60677678 -1.09817231 0 0 Z " fill="#DDE4E4" transform="translate(568,724)"/>
<path d="M0 0 C2.475 0.99 2.475 0.99 5 2 C2.42033404 4.57966596 -0.09307892 5.33609844 -3.5 6.625 C-4.6653125 7.07101562 -5.830625 7.51703125 -7.03125 7.9765625 C-10 9 -10 9 -12 9 C-11.34 7.02 -10.68 5.04 -10 3 C-8.3603125 3.0928125 -8.3603125 3.0928125 -6.6875 3.1875 C-3.07873917 3.35597914 -3.07873917 3.35597914 -1.0625 1.5 C-0.711875 1.005 -0.36125 0.51 0 0 Z " fill="#D5DDDD" transform="translate(604,696)"/>
<path d="M0 0 C5.67865696 2.47531201 10.20732567 6.1126086 15 10 C14.67 11.32 14.34 12.64 14 14 C13.01 14 12.02 14 11 14 C10.67 12.35 10.34 10.7 10 9 C9.01 9 8.02 9 7 9 C6.67 8.34 6.34 7.68 6 7 C5.360625 6.9175 4.72125 6.835 4.0625 6.75 C3.381875 6.5025 2.70125 6.255 2 6 C0.75 2.9375 0.75 2.9375 0 0 Z " fill="#D34B79" transform="translate(629,298)"/>
<path d="M0 0 C4.29 0.99 8.58 1.98 13 3 C9.41090147 5.39273235 7.73686522 6.15310986 3.5 6.1875 C2.7059375 6.20167969 1.911875 6.21585938 1.09375 6.23046875 C-1 6 -1 6 -3 4 C-2.01 2.68 -1.02 1.36 0 0 Z " fill="#DEE5E4" transform="translate(569,242)"/>
<path d="M0 0 C0 3.60777515 -0.9904432 5.06295544 -3 8 C-3.99 8.495 -3.99 8.495 -5 9 C-5 9.99 -5 10.98 -5 12 C-5.66 12 -6.32 12 -7 12 C-7.66 13.32 -8.32 14.64 -9 16 C-9.99 15.67 -10.98 15.34 -12 15 C-12.99 15 -13.98 15 -15 15 C-10.05 10.05 -5.1 5.1 0 0 Z " fill="#A32D6A" transform="translate(505,603)"/>
<path d="M0 0 C-1.43474844 4.09501116 -3.43465486 7.2603761 -6 10.75 C-6.70125 11.71421875 -7.4025 12.6784375 -8.125 13.671875 C-10 16 -10 16 -12 17 C-12.375 13.75 -12.375 13.75 -12 10 C-7.28205128 6 -7.28205128 6 -4 6 C-4 5.34 -4 4.68 -4 4 C-4.66 3.67 -5.32 3.34 -6 3 C-2.25 0 -2.25 0 0 0 Z " fill="#D46F96" transform="translate(701,583)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C-3.94 6.94 -9.88 12.88 -16 19 C-16.66 18.67 -17.32 18.34 -18 18 C-6.66287016 5.33029613 -6.66287016 5.33029613 0 0 Z " fill="#43C3A9" transform="translate(361,323)"/>
<path d="M0 0 C3.11601683 3.68256534 5.5162638 7.44792284 7.8125 11.6875 C8.43769531 12.82574219 9.06289063 13.96398437 9.70703125 15.13671875 C10.13371094 16.08160156 10.56039062 17.02648437 11 18 C10.67 18.66 10.34 19.32 10 20 C9.01 20 8.02 20 7 20 C6.87625 18.906875 6.7525 17.81375 6.625 16.6875 C6.24535199 12.92618198 6.24535199 12.92618198 4 10 C2.68 9.67 1.36 9.34 0 9 C0 6.03 0 3.06 0 0 Z " fill="#D3547B" transform="translate(689,358)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C3.19294408 5.82360189 2.75747614 9.49646738 1 14 C-0.96301592 10.49461443 -1.95902388 6.86648272 -3 3 C-2.01 2.01 -1.02 1.02 0 0 Z " fill="#CF5E87" transform="translate(729,498)"/>
<path d="M0 0 C0 3.26229641 -0.21770324 4.32655486 -2 7 C-3.3303125 7.86044922 -3.3303125 7.86044922 -4.6875 8.73828125 C-8.38536135 11.13215991 -11.32098776 14.09795774 -14.375 17.25 C-14.92027344 17.80429687 -15.46554687 18.35859375 -16.02734375 18.9296875 C-17.35622977 20.28188731 -18.67878548 21.6403035 -20 23 C-20.66 22.67 -21.32 22.34 -22 22 C-14.74 14.74 -7.48 7.48 0 0 Z " fill="#755892" transform="translate(320,460)"/>
<path d="M0 0 C0 3.77110589 -1.13327343 4.9680326 -3.3125 8 C-3.92738281 8.86625 -4.54226563 9.7325 -5.17578125 10.625 C-6.68648007 12.59181988 -8.19346467 14.31019465 -10 16 C-11.07425647 12.77723058 -11.26658842 12.03981221 -10 9 C-7.71484375 6.640625 -7.71484375 6.640625 -4.9375 4.25 C-4.01839844 3.45078125 -3.09929688 2.6515625 -2.15234375 1.828125 C-1.44207031 1.22484375 -0.73179687 0.6215625 0 0 Z " fill="#AA3969" transform="translate(716,511)"/>
<path d="M0 0 C3.63 0 7.26 0 11 0 C11.33 0.99 11.66 1.98 12 3 C11.67 3.66 11.34 4.32 11 5 C9.56208484 4.85831863 8.1246763 4.71148957 6.6875 4.5625 C5.88699219 4.48128906 5.08648437 4.40007813 4.26171875 4.31640625 C2 4 2 4 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#944C7D" transform="translate(448,680)"/>
<path d="M0 0 C2.66666667 2.66666667 5.33333333 5.33333333 8 8 C7.67 8.99 7.34 9.98 7 11 C2.93184627 9.15083921 -0.0094833 7.33557632 -3 4 C-2.34 4 -1.68 4 -1 4 C-0.67 2.68 -0.34 1.36 0 0 Z " fill="#763467" transform="translate(456,660)"/>
<path d="M0 0 C2 3 2 3 1.625 5.1875 C1.41875 5.785625 1.2125 6.38375 1 7 C-0.60875 7.37125 -0.60875 7.37125 -2.25 7.75 C-5.99649437 8.99883146 -7.52073882 10.02488658 -10 13 C-10.66 12.67 -11.32 12.34 -12 12 C-8.04 8.04 -4.08 4.08 0 0 Z " fill="#E3EAE8" transform="translate(700,646)"/>
<path d="M0 0 C1.16959987 0.97566112 2.33561177 1.955625 3.5 2.9375 C4.1496875 3.48277344 4.799375 4.02804687 5.46875 4.58984375 C6.22671875 5.28787109 6.22671875 5.28787109 7 6 C7 6.33 7 6.66 7 7 C5.8553125 6.938125 5.8553125 6.938125 4.6875 6.875 C1.77281584 6.77919176 1.77281584 6.77919176 -1 9 C-1 8.34 -1 7.68 -1 7 C-1.66 7 -2.32 7 -3 7 C-2.625 4.0625 -2.625 4.0625 -2 1 C-1.34 0.67 -0.68 0.34 0 0 Z " fill="#F2E4E9" transform="translate(648,488)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C-0.57871821 5.20430375 -2.14761637 7.16942403 -3.9375 9.1875 C-4.41896484 9.74630859 -4.90042969 10.30511719 -5.39648438 10.88085938 C-6.58857598 12.26179717 -7.79314375 13.63194679 -9 15 C-9.66 14.34 -10.32 13.68 -11 13 C-7.61227103 8.30840284 -4.21814817 3.9700218 0 0 Z " fill="#E2F8F5" transform="translate(338,344)"/>
<path d="M0 0 C0.99 0.66 1.98 1.32 3 2 C1.13133238 2.70453003 -0.74531416 3.38791688 -2.625 4.0625 C-3.66914062 4.44535156 -4.71328125 4.82820312 -5.7890625 5.22265625 C-9.30427743 6.07366327 -11.53329434 5.97088091 -15 5 C-15.33 4.34 -15.66 3.68 -16 3 C-14.39318359 2.80083984 -14.39318359 2.80083984 -12.75390625 2.59765625 C-11.35674231 2.4194944 -9.95960841 2.24109681 -8.5625 2.0625 C-7.85544922 1.97548828 -7.14839844 1.88847656 -6.41992188 1.79882812 C-2.91182032 1.61783809 -2.91182032 1.61783809 0 0 Z " fill="#D57497" transform="translate(590,670)"/>
<path d="M0 0 C0 3.10551666 -0.5393715 4.35261084 -2 7 C-2.66 7 -3.32 7 -4 7 C-4.33 7.99 -4.66 8.98 -5 10 C-7.875 12.25 -7.875 12.25 -11 14 C-11.99 13.67 -12.98 13.34 -14 13 C-9.38 8.71 -4.76 4.42 0 0 Z " fill="#215E59" transform="translate(683,648)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C-2.82320557 4.42258812 -5.91281305 5.24042276 -10 5 C-10 4.34 -10 3.68 -10 3 C-10.99 2.67 -11.98 2.34 -13 2 C-11.35524035 0.35524035 -9.32160131 0.64169424 -7.0625 0.4375 C-5.71865234 0.31181641 -5.71865234 0.31181641 -4.34765625 0.18359375 C-2 0 -2 0 0 0 Z " fill="#1B936E" transform="translate(476,343)"/>
<path d="M0 0 C0 3 0 3 -1 6 C-2.96317377 7.96317377 -4.61756195 9.57053717 -7 11 C-9.75 10.6875 -9.75 10.6875 -12 10 C-8.29909479 6.0747975 -4.45040344 3.05419844 0 0 Z " fill="#DCE3E1" transform="translate(374,276)"/>
<path d="M0 0 C1.32 0.33 2.64 0.66 4 1 C2.35 5.29 0.7 9.58 -1 14 C-1.66 13.01 -2.32 12.02 -3 11 C-2.125 8.3125 -2.125 8.3125 -1 6 C-1.66 6 -2.32 6 -3 6 C-3 5.01 -3 4.02 -3 3 C-2.34 3 -1.68 3 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#CFD9D5" transform="translate(739,556)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.85298376 3.67387495 2.10789471 7.0447393 2.0625 10.8125 C2.05347656 11.78832031 2.04445313 12.76414062 2.03515625 13.76953125 C2.02355469 14.50558594 2.01195312 15.24164063 2 16 C0.02 16.99 0.02 16.99 -2 18 C-1.48758893 11.97099313 -0.930215 5.97995357 0 0 Z " fill="#2D6662" transform="translate(259,430)"/>
<path d="M0 0 C2.31 0 4.62 0 7 0 C7.22174933 1.45635371 7.42698698 2.91522956 7.625 4.375 C7.74101563 5.18710937 7.85703125 5.99921875 7.9765625 6.8359375 C7.98429688 7.55007813 7.99203125 8.26421875 8 9 C7.34 9.66 6.68 10.32 6 11 C4.9944239 9.54550599 3.99569565 8.08627557 3 6.625 C2.443125 5.81289063 1.88625 5.00078125 1.3125 4.1640625 C0 2 0 2 0 0 Z " fill="#A72E69" transform="translate(617,392)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1 7.59 1 15.18 1 23 C0.67 23 0.34 23 0 23 C-0.13277344 21.99839844 -0.26554688 20.99679687 -0.40234375 19.96484375 C-0.58071127 18.62239346 -0.7590977 17.27994567 -0.9375 15.9375 C-1.02451172 15.28072266 -1.11152344 14.62394531 -1.20117188 13.94726562 C-1.77569697 9.62768808 -2.37745827 5.31292423 -3 1 C-2.01 1.33 -1.02 1.66 0 2 C0 1.34 0 0.68 0 0 Z " fill="#A42762" transform="translate(575,302)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.02724423 2.83339965 1.04695589 5.66653117 1.0625 8.5 C1.07087891 9.29148437 1.07925781 10.08296875 1.08789062 10.8984375 C1.10891185 16.02761717 0.73937287 20.92336106 0 26 C-1.64956143 23.03078942 -2.66052758 20.39472417 -3 17 C-2.68804688 16.42765625 -2.37609375 15.8553125 -2.0546875 15.265625 C-0.64935589 12.2467645 -0.5737869 9.56311508 -0.375 6.25 C-0.30023437 5.07953125 -0.22546875 3.9090625 -0.1484375 2.703125 C-0.09945312 1.81109375 -0.05046875 0.9190625 0 0 Z " fill="#CDDDD8" transform="translate(755,481)"/>
<path d="M0 0 C1.125 3.75 1.125 3.75 0 6 C0.66 6 1.32 6 2 6 C1 8 0 10 -1 12 C-0.34 12.33 0.32 12.66 1 13 C-2 17.5 -2 17.5 -5 22 C-4.36684209 16.87475334 -3.31839344 12.03469229 -1.9375 7.0625 C-1.75123047 6.37865234 -1.56496094 5.69480469 -1.37304688 4.99023438 C-0.91910943 3.32579707 -0.46009084 1.66274688 0 0 Z " fill="#50CEB1" transform="translate(298,418)"/>
<path d="M0 0 C0.33 0.66 0.66 1.32 1 2 C0.22265625 3.7265625 0.22265625 3.7265625 -0.9375 5.625 C-1.618125 6.73875 -2.29875 7.8525 -3 9 C-2.34 9 -1.68 9 -1 9 C-1 9.99 -1 10.98 -1 12 C-2.98 12.66 -4.96 13.32 -7 14 C-7.66 13.34 -8.32 12.68 -9 12 C-6.03 8.04 -3.06 4.08 0 0 Z " fill="#3CC6A6" transform="translate(336,349)"/>
<path d="M0 0 C2.31 0 4.62 0 7 0 C7.33 1.32 7.66 2.64 8 4 C9.65 4 11.3 4 13 4 C13.33 5.65 13.66 7.3 14 9 C12.22566188 8.06915029 10.45564851 7.13005387 8.6875 6.1875 C7.70136719 5.66542969 6.71523438 5.14335938 5.69921875 4.60546875 C3.38334932 3.2280124 1.76388999 2.00469409 0 0 Z " fill="#CED9D8" transform="translate(375,678)"/>
<path d="M0 0 C3.15204981 1.39347376 5.26171773 3.02485079 7.671875 5.4765625 C8.33574219 6.146875 8.99960937 6.8171875 9.68359375 7.5078125 C10.36550781 8.20648438 11.04742187 8.90515625 11.75 9.625 C12.44738281 10.33140625 13.14476562 11.0378125 13.86328125 11.765625 C15.58012488 13.50598703 17.29211832 15.25084981 19 17 C14.09452071 17 11.38197584 13.30917402 8 10 C7.04193199 8.89246358 6.10130053 7.7693338 5.1875 6.625 C3.20286584 3.77520272 3.20286584 3.77520272 0 3 C0 2.01 0 1.02 0 0 Z " fill="#572E68" transform="translate(352,445)"/>
<path d="M0 0 C3.63559661 3.43361902 6.36113346 6.7973607 9 11 C7.125 11.625 7.125 11.625 5 12 C4.34 11.34 3.68 10.68 3 10 C3 8.68 3 7.36 3 6 C2.01 6 1.02 6 0 6 C0 4.02 0 2.04 0 0 Z " fill="#D5527C" transform="translate(674,338)"/>
<path d="M0 0 C0 0.99 0 1.98 0 3 C-0.5775 3.061875 -1.155 3.12375 -1.75 3.1875 C-4.26157843 3.84640764 -4.26157843 3.84640764 -5.75 6.5625 C-8 9 -8 9 -10.03125 9.328125 C-12.02378804 9.31409304 -14.01429543 9.16547538 -16 9 C-11.97806144 5.49702126 -5.60566856 0 0 0 Z " fill="#255A5A" transform="translate(394,253)"/>
<path d="M0 0 C2.1519437 3.22791555 2.20086443 4.28400809 2 8 C3.32 8.66 4.64 9.32 6 10 C5.01 10.66 4.02 11.32 3 12 C1.99406757 10.8803014 0.9954151 9.7540588 0 8.625 C-0.556875 7.99851562 -1.11375 7.37203125 -1.6875 6.7265625 C-3 5 -3 5 -3 3 C-2.34 3 -1.68 3 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#D7719A" transform="translate(478,643)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C-0.8125 5.6875 -0.8125 5.6875 -3 8 C-3.66 8 -4.32 8 -5 8 C-6.59108002 9.44748074 -8.12559489 10.95775474 -9.625 12.5 C-10.44226563 13.3353125 -11.25953125 14.170625 -12.1015625 15.03125 C-12.72804688 15.6809375 -13.35453125 16.330625 -14 17 C-14.66 16.67 -15.32 16.34 -16 16 C-10.72 10.72 -5.44 5.44 0 0 Z " fill="#CBD9D7" transform="translate(343,301)"/>
<path d="M0 0 C2.31 0.33 4.62 0.66 7 1 C9.125 5.625 9.125 5.625 8 9 C5.03 7.02 2.06 5.04 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#A8356D" transform="translate(582,359)"/>
<path d="M0 0 C1.65 0.33 3.3 0.66 5 1 C-0.0022779 11.74259681 -0.0022779 11.74259681 -4 15 C-2.24215247 8.47085202 -2.24215247 8.47085202 -0.875 5.8125 C0.28983271 3.73507479 0.28983271 3.73507479 0 0 Z " fill="#D36F96" transform="translate(705,568)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C2.67 2.65 2.34 4.3 2 6 C1.01 6.33 0.02 6.66 -1 7 C-1.66 7.99 -2.32 8.98 -3 10 C-3.75 7.8125 -3.75 7.8125 -4 5 C-2.0625 2.1875 -2.0625 2.1875 0 0 Z " fill="#A62B64" transform="translate(629,547)"/>
<path d="M0 0 C-0.33 1.65 -0.66 3.3 -1 5 C-1.33 4.34 -1.66 3.68 -2 3 C-2.68707031 3.09539062 -3.37414062 3.19078125 -4.08203125 3.2890625 C-4.98308594 3.39992188 -5.88414062 3.51078125 -6.8125 3.625 C-7.70582031 3.74101562 -8.59914063 3.85703125 -9.51953125 3.9765625 C-12 4 -12 4 -15 2 C-13.43883181 1.66048381 -11.87598662 1.32867456 -10.3125 1 C-9.44238281 0.814375 -8.57226562 0.62875 -7.67578125 0.4375 C-5.06287036 0.01027953 -2.64186962 -0.07616201 0 0 Z " fill="#E4F7F3" transform="translate(486,345)"/>
<path d="M0 0 C2.3125 1.3125 2.3125 1.3125 3.3125 4.3125 C4.3025 4.3125 5.2925 4.3125 6.3125 4.3125 C6.3125 4.9725 6.3125 5.6325 6.3125 6.3125 C1.45286821 5.70504603 -2.4280518 3.58491033 -6.6875 1.3125 C-3.0234375 -0.7734375 -3.0234375 -0.7734375 0 0 Z " fill="#CAD6D5" transform="translate(399.6875,688.6875)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C2.61479436 3.53910197 2.29902057 4.72751123 0.37109375 6.484375 C-0.26699219 6.90203125 -0.90507812 7.3196875 -1.5625 7.75 C-2.20316406 8.17796875 -2.84382813 8.6059375 -3.50390625 9.046875 C-4.24447266 9.51867187 -4.24447266 9.51867187 -5 10 C-5.66 9.67 -6.32 9.34 -7 9 C-4.69 6.03 -2.38 3.06 0 0 Z " fill="#CFDAD9" transform="translate(314,334)"/>
<path d="M0 0 C0.33 0.66 0.66 1.32 1 2 C1.66 2.33 2.32 2.66 3 3 C2.40844669 4.31823302 1.80128537 5.62947051 1.1875 6.9375 C0.85105469 7.66839844 0.51460938 8.39929688 0.16796875 9.15234375 C-1 11 -1 11 -4 12 C-3.33501617 7.61110675 -1.81242323 4.0188515 0 0 Z " fill="#255854" transform="translate(276,377)"/>
<path d="M0 0 C0 3 0 3 -2.3125 5.625 C-5 8 -5 8 -8 9 C-8.33 9.66 -8.66 10.32 -9 11 C-9.99 10.67 -10.98 10.34 -12 10 C-8.04 6.7 -4.08 3.4 0 0 Z " fill="#48C6A8" transform="translate(376,310)"/>
<path d="M0 0 C2.31 0 4.62 0 7 0 C6.42655063 2.86724686 6.1385485 3.8614515 4 6 C1.525 5.01 1.525 5.01 -1 4 C-0.67 2.68 -0.34 1.36 0 0 Z " fill="#E9F0F0" transform="translate(609,240)"/>
<path d="M0 0 C1.55053541 4.65160624 1.82489894 9.93775265 0 14.5 C-0.33 14.995 -0.66 15.49 -1 16 C-3.48824257 12.26763615 -2.99011601 11.1728793 -2.1875 6.875 C-1.99542969 5.79992187 -1.80335938 4.72484375 -1.60546875 3.6171875 C-1 1 -1 1 0 0 Z " fill="#D36490" transform="translate(722,528)"/>
<path d="M0 0 C1.67110042 2.96178773 2.32682752 5.37071192 2.625 8.75 C2.69976563 9.54921875 2.77453125 10.3484375 2.8515625 11.171875 C2.90054688 11.77515625 2.94953125 12.3784375 3 13 C1.68 12.67 0.36 12.34 -1 12 C-1.14285714 3.42857143 -1.14285714 3.42857143 0 0 Z " fill="#DC6187" transform="translate(715,417)"/>
<path d="M0 0 C0 2.64 0 5.28 0 8 C-1.17219543 7.21654285 -2.33763668 6.42297164 -3.5 5.625 C-4.1496875 5.18414062 -4.799375 4.74328125 -5.46875 4.2890625 C-5.9740625 3.86367188 -6.479375 3.43828125 -7 3 C-7 2.34 -7 1.68 -7 1 C-4 0 -4 0 0 0 Z " fill="#A12C65" transform="translate(601,368)"/>
<path d="M0 0 C3.3 0 6.6 0 10 0 C9 2 9 2 6.75 3.1875 C3.69751418 4.08937081 2.02265546 3.86361585 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#D1DAD9" transform="translate(575,706)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C2.49477778 5.37859255 -0.17827222 7.81651224 -3 11 C-4 8 -4 8 -3.22265625 5.95703125 C-2.83980469 5.24933594 -2.45695313 4.54164063 -2.0625 3.8125 C-1.68222656 3.09707031 -1.30195312 2.38164063 -0.91015625 1.64453125 C-0.60980469 1.10183594 -0.30945313 0.55914063 0 0 Z " fill="#A63B6A" transform="translate(641,523)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C-0.63 4.3 -4.26 7.6 -8 11 C-8.33 10.01 -8.66 9.02 -9 8 C-8.34 8 -7.68 8 -7 8 C-6.67 7.01 -6.34 6.02 -6 5 C-3.125 2.25 -3.125 2.25 0 0 Z " fill="#D65A83" transform="translate(696,496)"/>
<path d="M0 0 C1.65 0.33 3.3 0.66 5 1 C4.01 2.98 3.02 4.96 2 7 C-0.97 6.505 -0.97 6.505 -4 6 C-3.34 5.67 -2.68 5.34 -2 5 C-1.27840576 3.35636866 -0.60648579 1.68949614 0 0 Z " fill="#E3EBE9" transform="translate(595,232)"/>
<path d="M0 0 C0.33 0.66 0.66 1.32 1 2 C3.02463255 2.65213292 3.02463255 2.65213292 5 3 C3.71086513 3.67154933 2.41859796 4.33708859 1.125 5 C0.40570312 5.37125 -0.31359375 5.7425 -1.0546875 6.125 C-3 7 -3 7 -5 7 C-4.75 4.625 -4.75 4.625 -4 2 C-1.9375 0.6875 -1.9375 0.6875 0 0 Z " fill="#CED8D7" transform="translate(621,688)"/>
<path d="M0 0 C2.56616632 3.84924948 2.55097676 6.4349304 3 11 C2.01 11 1.02 11 0 11 C-1.76062164 7.67438135 -2.10784228 6.40826005 -1.125 2.6875 C-0.568125 1.3571875 -0.568125 1.3571875 0 0 Z " fill="#2D6866" transform="translate(756,406)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C0.71937515 2.7074998 -0.61767557 4.37373596 -2 6 C-2.66 6 -3.32 6 -4 6 C-4 6.66 -4 7.32 -4 8 C-5.65 7.67 -7.3 7.34 -9 7 C-6.03716687 4.61327331 -3.05729491 2.2646629 0 0 Z " fill="#45C6A3" transform="translate(389,301)"/>
<path d="M0 0 C1.98 0.99 3.96 1.98 6 3 C5.67 4.32 5.34 5.64 5 7 C3.35 6.67 1.7 6.34 0 6 C0 4.02 0 2.04 0 0 Z " fill="#A52E64" transform="translate(648,529)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C2.01 4.96 1.02 8.92 0 13 C-2.0903754 8.81924919 -2.22667078 8.41186737 -1.125 4.25 C-0.92132812 3.45078125 -0.71765625 2.6515625 -0.5078125 1.828125 C-0.34023438 1.22484375 -0.17265625 0.6215625 0 0 Z " fill="#D7749B" transform="translate(724,524)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C1.34 2.31 0.68 4.62 0 7 C-3 7 -3 7 -5.1875 5.125 C-7 3 -7 3 -7 1 C-6.34 1 -5.68 1 -5 1 C-5 1.66 -5 2.32 -5 3 C-3.02463255 2.65213292 -3.02463255 2.65213292 -1 2 C-0.67 1.34 -0.34 0.68 0 0 Z " fill="#219F86" transform="translate(382,423)"/>
<path d="M0 0 C0.66 0.66 1.32 1.32 2 2 C0.92319498 3.13125022 -0.16175635 4.25474919 -1.25 5.375 C-1.85328125 6.00148438 -2.4565625 6.62796875 -3.078125 7.2734375 C-4.9700588 8.97310161 -6.68201309 9.98459866 -9 11 C-8.46324097 7.14896699 -6.88399077 5.68202413 -3.9375 3.25 C-3.20402344 2.63640625 -2.47054688 2.0228125 -1.71484375 1.390625 C-1.14894531 0.93171875 -0.58304687 0.4728125 0 0 Z " fill="#DBF6F3" transform="translate(366,315)"/>
<path d="M0 0 C2.475 0.99 2.475 0.99 5 2 C5 2.99 5 3.98 5 5 C6.32 5.66 7.64 6.32 9 7 C9 7.99 9 8.98 9 10 C4.50486731 8.50162244 2.37078067 4.87680938 0 1 C0 0.67 0 0.34 0 0 Z " fill="#D2DCDC" transform="translate(312,618)"/>
<path d="M0 0 C2.475 0.99 2.475 0.99 5 2 C4.67 4.64 4.34 7.28 4 10 C1.7448078 7.7448078 1.02276532 5.9952413 0 3 C0 2.01 0 1.02 0 0 Z " fill="#D4DDDD" transform="translate(281,561)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C2.20568053 4.67201205 2.09382426 9.21496292 2 14 C1.01 13.67 0.02 13.34 -1 13 C-0.67 8.71 -0.34 4.42 0 0 Z " fill="#1F5F59" transform="translate(755,499)"/>
<path d="M0 0 C0.66 0.66 1.32 1.32 2 2 C-1.96 3.98 -1.96 3.98 -6 6 C-6.99 5.34 -7.98 4.68 -9 4 C-8.34 4 -7.68 4 -7 4 C-7 3.34 -7 2.68 -7 2 C-4.69 1.34 -2.38 0.68 0 0 Z " fill="#E1ECED" transform="translate(372,263)"/>
<path d="M0 0 C1 2 1 2 0.3125 4.5 C-1 7 -1 7 -2.9375 8.375 C-5 9 -5 9 -8 8 C-5.36 5.36 -2.72 2.72 0 0 Z " fill="#A63470" transform="translate(489,619)"/>
<path d="M0 0 C1.32 0 2.64 0 4 0 C4.33 0.99 4.66 1.98 5 3 C5.66 3.66 6.32 4.32 7 5 C4.69 5.33 2.38 5.66 0 6 C0 4.02 0 2.04 0 0 Z " fill="#EBE3E7" transform="translate(536,601)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C-1.25 4.625 -1.25 4.625 -4 6 C-6.3125 5.1875 -6.3125 5.1875 -8 4 C-3.375 0 -3.375 0 0 0 Z " fill="#E2EDEB" transform="translate(393,250)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C1.71372289 2.17260611 0.42080217 3.3379283 -0.875 4.5 C-1.59429688 5.1496875 -2.31359375 5.799375 -3.0546875 6.46875 C-5 8 -5 8 -7 8 C-5.51218185 4.21282653 -3.38011591 2.22592999 0 0 Z " fill="#9D2860" transform="translate(704,522)"/>
<path d="M0 0 C1.0625 1.875 1.0625 1.875 2 4 C1.67 4.66 1.34 5.32 1 6 C0.34 6 -0.32 6 -1 6 C-1.66 7.98 -2.32 9.96 -3 12 C-3.66 12 -4.32 12 -5 12 C-3.68938409 7.76570244 -2.05643741 3.92592596 0 0 Z " fill="#54CAB0" transform="translate(312,385)"/>
<path d="M0 0 C1.65 0 3.3 0 5 0 C5 2.31 5 4.62 5 7 C3.02 5.35 1.04 3.7 -1 2 C-0.67 1.34 -0.34 0.68 0 0 Z " fill="#9E235E" transform="translate(604,376)"/>
<path d="M0 0 C0.99 0.66 1.98 1.32 3 2 C2.01 2.495 2.01 2.495 1 3 C1 4.32 1 5.64 1 7 C-0.98 7.99 -0.98 7.99 -3 9 C-3.75 6.75 -3.75 6.75 -4 4 C-2.0625 1.6875 -2.0625 1.6875 0 0 Z " fill="#1B5854" transform="translate(285,362)"/>
<path d="M0 0 C0 0.99 0 1.98 0 3 C-0.639375 3.268125 -1.27875 3.53625 -1.9375 3.8125 C-4.33131686 4.88667752 -4.33131686 4.88667752 -5 8 C-6.65 8.33 -8.3 8.66 -10 9 C-6.83047153 5.73991357 -3.60062011 2.77762123 0 0 Z " fill="#285959" transform="translate(354,278)"/>
<path d="M0 0 C0.66 1.32 1.32 2.64 2 4 C2.66 4.33 3.32 4.66 4 5 C3.67 6.98 3.34 8.96 3 11 C2.01 11 1.02 11 0 11 C0 7.37 0 3.74 0 0 Z " fill="#3AC38F" transform="translate(484,260)"/>
<path d="M0 0 C1.98 0 3.96 0 6 0 C6 0.99 6 1.98 6 3 C5.01 3 4.02 3 3 3 C3 3.66 3 4.32 3 5 C1.68 4.67 0.36 4.34 -1 4 C-0.67 2.68 -0.34 1.36 0 0 Z " fill="#EAF2F3" transform="translate(626,248)"/>
<path d="M0 0 C0 0.33 0 0.66 0 1 C-3.96 1.66 -7.92 2.32 -12 3 C-12 2.01 -12 1.02 -12 0 C-7.6835078 -0.76173392 -4.25566547 -1.16063604 0 0 Z " fill="#DFEFED" transform="translate(464,228)"/>
<path d="M0 0 C2.96175123 0.61277612 4.38058783 1.25372522 7 3 C6 4 6 4 3.93359375 4.09765625 C3.10988281 4.08605469 2.28617188 4.07445312 1.4375 4.0625 C0.61121094 4.05347656 -0.21507812 4.04445313 -1.06640625 4.03515625 C-1.70449219 4.02355469 -2.34257813 4.01195312 -3 4 C-2.67 3.34 -2.34 2.68 -2 2 C-1.34 2 -0.68 2 0 2 C0 1.34 0 0.68 0 0 Z " fill="#A52A63" transform="translate(549,604)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.05416188 1.60379341 1.09286638 3.20811406 1.125 4.8125 C1.14820313 5.70582031 1.17140625 6.59914063 1.1953125 7.51953125 C1 10 1 10 -1 13 C-1.66 13 -2.32 13 -3 13 C-2.01 8.71 -1.02 4.42 0 0 Z " fill="#D0DEDC" transform="translate(277,403)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C2 0.66 2 1.32 2 2 C3.32 1.67 4.64 1.34 6 1 C6 2.65 6 4.3 6 6 C5.01 6.33 4.02 6.66 3 7 C0 2.25 0 2.25 0 0 Z " fill="#A32663" transform="translate(626,405)"/>
<path d="M0 0 C2.22825644 2.22825644 2.69239369 3.65761628 3.625 6.625 C4.01558594 7.85089844 4.01558594 7.85089844 4.4140625 9.1015625 C4.60742188 9.72804688 4.80078125 10.35453125 5 11 C4.01 11 3.02 11 2 11 C0.80712589 7.12315913 0 4.08378077 0 0 Z " fill="#D35980" transform="translate(703,384)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C0.78192862 2.15762119 -0.45001235 3.3006583 -1.6875 4.4375 C-2.71423828 5.39462891 -2.71423828 5.39462891 -3.76171875 6.37109375 C-6.22289422 8.16221098 -8.00816574 8.62798558 -11 9 C-7.56638098 5.36440339 -4.2026393 2.63886654 0 0 Z " fill="#CFF0EA" transform="translate(437,362)"/>
<path d="M0 0 C0.33 1.32 0.66 2.64 1 4 C0.01 4 -0.98 4 -2 4 C-4.17032476 5.43990623 -4.17032476 5.43990623 -6 7 C-7.32 6.34 -8.64 5.68 -10 5 C-6.7 3.35 -3.4 1.7 0 0 Z " fill="#D2DCDC" transform="translate(402,260)"/>
<path d="M0 0 C2.02054804 1.64169528 4.02043058 3.30911778 6 5 C6 5.33 6 5.66 6 6 C3.03 6 0.06 6 -3 6 C-2.01 5.67 -1.02 5.34 0 5 C-0.2784375 4.0409375 -0.2784375 4.0409375 -0.5625 3.0625 C-0.706875 2.381875 -0.85125 1.70125 -1 1 C-0.67 0.67 -0.34 0.34 0 0 Z " fill="#A0E6CF" transform="translate(495,253)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.125 2.375 1.125 2.375 1 5 C0.34 5.66 -0.32 6.32 -1 7 C-3.625 6.625 -3.625 6.625 -6 6 C-4 3 -4 3 -1 2 C-0.67 1.34 -0.34 0.68 0 0 Z " fill="#D27E9A" transform="translate(536,699)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C0.515 3.475 0.515 3.475 -1 6 C-3.4375 5.625 -3.4375 5.625 -6 5 C-6.33 4.34 -6.66 3.68 -7 3 C-4.69631264 1.93347808 -2.35981813 0.93578995 0 0 Z " fill="#235C58" transform="translate(611,697)"/>
<path d="M0 0 C0 3.58912412 -0.66436554 4.10857029 -3 6.6875 C-3.556875 7.31011719 -4.11375 7.93273437 -4.6875 8.57421875 C-5.120625 9.04472656 -5.55375 9.51523437 -6 10 C-6.99 9.67 -7.98 9.34 -9 9 C-6.03 6.03 -3.06 3.06 0 0 Z " fill="#AA376D" transform="translate(615,564)"/>
<path d="M0 0 C1.9375 0.9375 1.9375 0.9375 4 3 C4.66174825 5.9858081 4.87205948 8.94861869 5 12 C1.94063363 8.24532309 0 4.91886939 0 0 Z " fill="#6D5289" transform="translate(316,560)"/>
<path d="M0 0 C2 2 2 2 2 6 C0.02 6.66 -1.96 7.32 -4 8 C-2.87548273 5.0280615 -1.77706209 2.66559313 0 0 Z " fill="#41CAA9" transform="translate(323,367)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C-0.75 7.875 -0.75 7.875 -3 9 C-3.66 8.67 -4.32 8.34 -5 8 C-3.8141763 4.62496331 -2.72426311 2.35277269 0 0 Z " fill="#A43D71" transform="translate(565,343)"/>
<path d="M0 0 C0.99 0 1.98 0 3 0 C3 0.66 3 1.32 3 2 C3.66 2 4.32 2 5 2 C6.625 4.5 6.625 4.5 8 7 C5 7 5 7 2.3125 4.625 C0 2 0 2 0 0 Z " fill="#C94F7C" transform="translate(546,272)"/>
<path d="M0 0 C0 0.99 0 1.98 0 3 C-2.64 3 -5.28 3 -8 3 C-8 2.34 -8 1.68 -8 1 C-3.375 -1.125 -3.375 -1.125 0 0 Z " fill="#8F5079" transform="translate(482,687)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C-1.3431213 2.74438677 -3.67843403 2.40729228 -6 2 C-6.33 1.34 -6.66 0.68 -7 0 C-3.89953913 -1.03348696 -2.94389782 -1.17755913 0 0 Z " fill="#864075" transform="translate(416,665)"/>
<path d="M0 0 C2.16874252 0.50603992 3.99967627 0.99983813 6 2 C5.67 3.98 5.34 5.96 5 8 C2.74754119 5.31158141 1.11786042 3.35358125 0 0 Z " fill="#D0DDDD" transform="translate(301,602)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C1.4409112 3.24271506 0.5867822 4.93057424 -2 7 C-2.66 7 -3.32 7 -4 7 C-4.33 7.66 -4.66 8.32 -5 9 C-4.38722388 6.03824877 -3.74627478 4.61941217 -2 2 C-1.34 2 -0.68 2 0 2 C0 1.34 0 0.68 0 0 Z " fill="#D95B86" transform="translate(739,453)"/>
<path d="M0 0 C2.05078125 0.03255208 4.1015625 0.06510417 6.15234375 0.09765625 C6.15234375 0.75765625 6.15234375 1.41765625 6.15234375 2.09765625 C2.77734375 2.72265625 2.77734375 2.72265625 -0.84765625 3.09765625 C-1.50765625 2.43765625 -2.16765625 1.77765625 -2.84765625 1.09765625 C-1.84765625 0.09765625 -1.84765625 0.09765625 0 0 Z " fill="#189470" transform="translate(447.84765625,351.90234375)"/>
<path d="M0 0 C0.66 0.66 1.32 1.32 2 2 C1.64644564 4.26274788 1.02455574 5.95088852 0 8 C-0.99 8 -1.98 8 -3 8 C-1.125 2.25 -1.125 2.25 0 0 Z " fill="#1E5C58" transform="translate(732,581)"/>
<path d="M0 0 C1.32 0.33 2.64 0.66 4 1 C3.01 2.32 2.02 3.64 1 5 C0.67 4.67 0.34 4.34 0 4 C-0.33 4.66 -0.66 5.32 -1 6 C-1.66 6 -2.32 6 -3 6 C-3 5.01 -3 4.02 -3 3 C-2.34 3 -1.68 3 -1 3 C-0.67 2.01 -0.34 1.02 0 0 Z " fill="#D9DFDD" transform="translate(739,556)"/>
<path d="M0 0 C1.65 0 3.3 0 5 0 C3.35 1.98 1.7 3.96 0 6 C-0.66 5.67 -1.32 5.34 -2 5 C-1.34 3.35 -0.68 1.7 0 0 Z " fill="#37B19A" transform="translate(311,434)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C2 0.66 2 1.32 2 2 C2.66 2 3.32 2 4 2 C4.625 4.8125 4.625 4.8125 5 8 C4.01 9.485 4.01 9.485 3 11 C2.01 7.37 1.02 3.74 0 0 Z " fill="#AB4176" transform="translate(634,422)"/>
<path d="M0 0 C-0.66 1.32 -1.32 2.64 -2 4 C-2.66 3.67 -3.32 3.34 -4 3 C-4.33 3.66 -4.66 4.32 -5 5 C-5.33 3.35 -5.66 1.7 -6 0 C-3.50907189 -1.24546405 -2.58919267 -0.7767578 0 0 Z " fill="#E4EAE9" transform="translate(296,340)"/>
<path d="M0 0 C0 0.66 0 1.32 0 2 C0.66 2 1.32 2 2 2 C2 2.66 2 3.32 2 4 C-2.455 3.01 -2.455 3.01 -7 2 C-4 0 -4 0 0 0 Z " fill="#CFD9DA" transform="translate(437,704)"/>
<path d="M0 0 C3.3 0 6.6 0 10 0 C8.68 0.33 7.36 0.66 6 1 C6 1.99 6 2.98 6 4 C4.68 3.67 3.36 3.34 2 3 C2 2.34 2 1.68 2 1 C1.34 0.67 0.68 0.34 0 0 Z " fill="#7B5E97" transform="translate(340,442)"/>
<path d="M0 0 C0.99 0.33 1.98 0.66 3 1 C2.01 3.97 1.02 6.94 0 10 C-0.66 10 -1.32 10 -2 10 C-1.34 6.7 -0.68 3.4 0 0 Z " fill="#C9D5D5" transform="translate(273,418)"/>
<path d="M0 0 C2.15377564 2.62198774 3.40072174 4.64404172 4 8 C3.01 8.33 2.02 8.66 1 9 C-1.125 2.25 -1.125 2.25 0 0 Z " fill="#C5D6D3" transform="translate(731,371)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C2.5625 3.3125 2.5625 3.3125 3 6 C3.32483418 7.33542939 3.6550855 8.66961551 4 10 C1.4375 7.8125 1.4375 7.8125 -1 5 C-0.8125 2.1875 -0.8125 2.1875 0 0 Z " fill="#A42D60" transform="translate(566,289)"/>
<path d="M0 0 C-0.66 1.32 -1.32 2.64 -2 4 C-2 3.34 -2 2.68 -2 2 C-2.7425 2.350625 -3.485 2.70125 -4.25 3.0625 C-7.21122875 4.0720098 -8.12062561 3.87980884 -11 3 C-9.73160474 2.49384702 -8.46016898 1.99530901 -7.1875 1.5 C-6.12595703 1.08234375 -6.12595703 1.08234375 -5.04296875 0.65625 C-3 0 -3 0 0 0 Z " fill="#B9CACB" transform="translate(438,246)"/>
<path d="M0 0 C1.9375 0.125 1.9375 0.125 4 1 C5.25 3.5625 5.25 3.5625 6 6 C5.01 6 4.02 6 3 6 C0.8125 3.5 0.8125 3.5 -1 1 C-0.67 0.67 -0.34 0.34 0 0 Z " fill="#DBE2E4" transform="translate(329,637)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.9765625 6.0546875 1.9765625 6.0546875 2 8 C1.34 8.66 0.68 9.32 0 10 C-1.49106457 7.01787087 -1.11941467 4.28390342 -1 1 C-0.67 0.67 -0.34 0.34 0 0 Z " fill="#E2EAE9" transform="translate(261,533)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C1.67 2.64 1.34 5.28 1 8 C0.01 6.68 -0.98 5.36 -2 4 C-1.34 2.68 -0.68 1.36 0 0 Z " fill="#D8E0DD" transform="translate(748,529)"/>
<path d="M0 0 C0.6875 1.6875 0.6875 1.6875 1 4 C-0.4375 6.75 -0.4375 6.75 -2 9 C-2.66 8.67 -3.32 8.34 -4 8 C-3.835 7.38125 -3.67 6.7625 -3.5 6.125 C-2.92365356 4.03936614 -2.92365356 4.03936614 -3 2 C-2.01 1.34 -1.02 0.68 0 0 Z " fill="#EDD7DC" transform="translate(489,421)"/>
<path d="M0 0 C0.66 0.66 1.32 1.32 2 2 C1.625 5.625 1.625 5.625 1 9 C-1 7 -1 7 -1.1875 3.9375 C-1 1 -1 1 0 0 Z " fill="#DAE3E1" transform="translate(260,417)"/>
<path d="M0 0 C1.65 1.65 3.3 3.3 5 5 C3.02 5.99 3.02 5.99 1 7 C0 6 0 6 -0.0625 2.9375 C-0.041875 1.968125 -0.02125 0.99875 0 0 Z " fill="#C7D6D4" transform="translate(710,337)"/>
<path d="M0 0 C0 0.99 0 1.98 0 3 C-2.25 4.75 -2.25 4.75 -5 6 C-6.32 5.67 -7.64 5.34 -9 5 C-6.03 3.35 -3.06 1.7 0 0 Z " fill="#4AC5A2" transform="translate(400,295)"/>
<path d="M0 0 C3 3.75 3 3.75 3 6 C4.32 6.33 5.64 6.66 7 7 C4.69 7 2.38 7 0 7 C0 4.69 0 2.38 0 0 Z " fill="#A4E2CC" transform="translate(484,252)"/>
<path d="M0 0 C2.31 0 4.62 0 7 0 C6.67 1.32 6.34 2.64 6 4 C3.69 3.34 1.38 2.68 -1 2 C-0.67 1.34 -0.34 0.68 0 0 Z " fill="#C5D2D1" transform="translate(423,701)"/>
<path d="M0 0 C1.98 0 3.96 0 6 0 C6 1.98 6 3.96 6 6 C3.97945196 4.35830472 1.97956942 2.69088222 0 1 C0 0.67 0 0.34 0 0 Z " fill="#D67497" transform="translate(505,678)"/>
<path d="M0 0 C0.33 0.99 0.66 1.98 1 3 C0.01 4.485 0.01 4.485 -1 6 C-3.625 6.1875 -3.625 6.1875 -6 6 C-4 4 -2 2 0 0 Z " fill="#B03F72" transform="translate(602,576)"/>
<path d="M0 0 C1.32 0.33 2.64 0.66 4 1 C3.34 2.98 2.68 4.96 2 7 C0 4 0 4 0 0 Z " fill="#6E528D" transform="translate(309,539)"/>
<path d="M0 0 C-1.39332574 3.36720387 -2.9789286 4.9859524 -6 7 C-5.37162381 3.35541809 -4.14650034 0 0 0 Z " fill="#D85A83" transform="translate(705,489)"/>
<path d="M0 0 C1.98 0 3.96 0 6 0 C6 0.99 6 1.98 6 3 C3.69 2.67 1.38 2.34 -1 2 C-0.67 1.34 -0.34 0.68 0 0 Z " fill="#F8F7F8" transform="translate(568,357)"/>
<path d="M0 0 C2.25 1.9375 2.25 1.9375 4 4 C-1.75 4.125 -1.75 4.125 -4 3 C-4 2.34 -4 1.68 -4 1 C-2.25 0.25 -2.25 0.25 0 0 Z " fill="#DEE7E4" transform="translate(668,292)"/>
<path d="M0 0 C0.66 0.33 1.32 0.66 2 1 C1.67 1.99 1.34 2.98 1 4 C-2.28976808 5.09658936 -3.71303767 4.79953138 -7 4 C-6.1028125 3.566875 -6.1028125 3.566875 -5.1875 3.125 C-2.80672208 1.95257974 -2.80672208 1.95257974 0 0 Z " fill="#31C394" transform="translate(432,283)"/>
<path d="M0 0 C0 0.99 0 1.98 0 3 C-2.3125 5.25 -2.3125 5.25 -5 7 C-5.99 6.67 -6.98 6.34 -8 6 C-5.36 4.02 -2.72 2.04 0 0 Z " fill="#CDDADA" transform="translate(374,276)"/>
<path d="M0 0 C-1.423125 0.680625 -1.423125 0.680625 -2.875 1.375 C-6.00313679 2.80238254 -6.00313679 2.80238254 -8 5 C-8.66 4.01 -9.32 3.02 -10 2 C-3.375 -1.125 -3.375 -1.125 0 0 Z " fill="#C9D7D8" transform="translate(427,251)"/>
<path d="M0 0 C-2.62198774 2.15377564 -4.64404172 3.40072174 -8 4 C-8.33 3.34 -8.66 2.68 -9 2 C-3.375 -1.125 -3.375 -1.125 0 0 Z " fill="#2B5D5B" transform="translate(403,250)"/>
<path d="M0 0 C2.33944736 0.28730055 4.6739143 0.61936779 7 1 C5.68 1.99 4.36 2.98 3 4 C1.68 3.01 0.36 2.02 -1 1 C-0.67 0.67 -0.34 0.34 0 0 Z " fill="#D7DEDE" transform="translate(631,682)"/>
<path d="M0 0 C2 2 2 2 2 5 C1.01 5.33 0.02 5.66 -1 6 C-1.99 4.68 -2.98 3.36 -4 2 C-3.34 1.67 -2.68 1.34 -2 1 C-1.34 1.33 -0.68 1.66 0 2 C0 1.34 0 0.68 0 0 Z " fill="#DFE5E4" transform="translate(344,648)"/>
<path d="M0 0 C0.33 0.66 0.66 1.32 1 2 C1.66 2 2.32 2 3 2 C2.34 4.97 1.68 7.94 1 11 C0.67 11 0.34 11 0 11 C0 7.37 0 3.74 0 0 Z " fill="#CE779F" transform="translate(474,635)"/>
<path d="M0 0 C2.475 0.99 2.475 0.99 5 2 C4.01 2.495 4.01 2.495 3 3 C3 3.66 3 4.32 3 5 C2.01 5 1.02 5 0 5 C0 3.35 0 1.7 0 0 Z " fill="#6A2662" transform="translate(432,586)"/>
<path d="M0 0 C0.66 0 1.32 0 2 0 C0.25 5.75 0.25 5.75 -2 8 C-3 5 -3 5 -1.6875 2.3125 C-1.130625 1.549375 -0.57375 0.78625 0 0 Z " fill="#CFDBD7" transform="translate(732,577)"/>
<path d="M0 0 C0.33 0 0.66 0 1 0 C1.125 3.375 1.125 3.375 1 7 C0.34 7.66 -0.32 8.32 -1 9 C-2.25541557 5.23375329 -1.37061958 3.62811066 0 0 Z " fill="#E4ECEB" transform="translate(264,404)"/>
<path d="M0 0 C-0.33 0.66 -0.66 1.32 -1 2 C-3.64 1.67 -6.28 1.34 -9 1 C-9 0.67 -9 0.34 -9 0 C-5.62182575 -0.84454356 -3.32534757 -1.10844919 0 0 Z " fill="#D7F3ED" transform="translate(480,347)"/>
<path d="M0 0 C0.99 0 1.98 0 3 0 C3.33 1.98 3.66 3.96 4 6 C2.02 5.01 0.04 4.02 -2 3 C-1.34 2.67 -0.68 2.34 0 2 C0 1.34 0 0.68 0 0 Z " fill="#DFE8E8" transform="translate(644,258)"/>
<path d="M0 0 C1.98 0.66 3.96 1.32 6 2 C4 4 4 4 1.375 4.125 C0.59125 4.08375 -0.1925 4.0425 -1 4 C-0.67 2.68 -0.34 1.36 0 0 Z " fill="#D2DADB" transform="translate(596,250)"/>
<path d="M0 0 C1.98 0 3.96 0 6 0 C5.67 1.32 5.34 2.64 5 4 C2.525 3.01 2.525 3.01 0 2 C0 1.34 0 0.68 0 0 Z " fill="#F6FBFB" transform="translate(407,240)"/>
<path d="M0 0 C-0.33 0.66 -0.66 1.32 -1 2 C-3.97 1.67 -6.94 1.34 -10 1 C-5.64467851 -1.17766075 -4.53374042 -1.03039555 0 0 Z " fill="#D5E3E2" transform="translate(570,229)"/>
</svg>
